// NIOS_Sys.v

// Generated using ACDS version 13.0sp1 232 at 2014.09.23.20:09:13

`timescale 1 ps / 1 ps
module NIOS_Sys (
		output wire [7:0]  led_external_connection_export,      //    led_external_connection.export
		output wire [12:0] sdram_wire_addr,                     //                 sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                       //                           .ba
		output wire        sdram_wire_cas_n,                    //                           .cas_n
		output wire        sdram_wire_cke,                      //                           .cke
		output wire        sdram_wire_cs_n,                     //                           .cs_n
		inout  wire [15:0] sdram_wire_dq,                       //                           .dq
		output wire [1:0]  sdram_wire_dqm,                      //                           .dqm
		output wire        sdram_wire_ras_n,                    //                           .ras_n
		output wire        sdram_wire_we_n,                     //                           .we_n
		input  wire [1:0]  key_external_connection_export,      //    key_external_connection.export
		input  wire [3:0]  sw_external_connection_export,       //     sw_external_connection.export
		input  wire        reset_reset_n,                       //                      reset.reset_n
		output wire        altpll_0_c1_clk,                     //                altpll_0_c1.clk
		input  wire        clk_clk,                             //                        clk.clk
		input  wire        ultrasound0_conduit_end_feedback_in, //    ultrasound0_conduit_end.feedback_in
		output wire        ultrasound0_conduit_end_trigger_out, //                           .trigger_out
		input  wire        ultrasound1_conduit_end_feedback_in, //    ultrasound1_conduit_end.feedback_in
		output wire        ultrasound1_conduit_end_trigger_out, //                           .trigger_out
		output wire        adc_spi_read_conduit_end_OUT,        //   adc_spi_read_conduit_end.OUT
		input  wire        adc_spi_read_conduit_end_IN,         //                           .IN
		output wire        adc_spi_read_conduit_end_CS_n,       //                           .CS_n
		output wire        adc_spi_read_conduit_end_CLK,        //                           .CLK
		output wire        pwm0_conduit_end_pwm1,               //           pwm0_conduit_end.pwm1
		output wire        pwm0_conduit_end_pwm2,               //                           .pwm2
		output wire        pwm1_conduit_end_pwm1,               //           pwm1_conduit_end.pwm1
		output wire        pwm1_conduit_end_pwm2,               //                           .pwm2
		input  wire [1:0]  encoder0_conduit_end_export,         //       encoder0_conduit_end.export
		input  wire [1:0]  encoder1_conduit_end_export,         //       encoder1_conduit_end.export
		output wire [7:0]  pio_0_external_connection_export,    //  pio_0_external_connection.export
		input  wire        uart_0_external_connection_rxd,      // uart_0_external_connection.rxd
		output wire        uart_0_external_connection_txd,      //                           .txd
		input  wire        ultrasound2_conduit_end_feedback_in, //    ultrasound2_conduit_end.feedback_in
		output wire        ultrasound2_conduit_end_trigger_out, //                           .trigger_out
		input  wire        ultrasound3_conduit_end_feedback_in, //    ultrasound3_conduit_end.feedback_in
		output wire        ultrasound3_conduit_end_trigger_out, //                           .trigger_out
		input  wire        ultrasound5_conduit_end_feedback_in, //    ultrasound5_conduit_end.feedback_in
		output wire        ultrasound5_conduit_end_trigger_out, //                           .trigger_out
		output wire        pwm2_conduit_end_pwm1,               //           pwm2_conduit_end.pwm1
		output wire        pwm2_conduit_end_pwm2,               //                           .pwm2
		output wire        pwm3_conduit_end_pwm1,               //           pwm3_conduit_end.pwm1
		output wire        pwm3_conduit_end_pwm2,               //                           .pwm2
		input  wire        ultrasound4_conduit_end_feedback_in, //    ultrasound4_conduit_end.feedback_in
		output wire        ultrasound4_conduit_end_trigger_out, //                           .trigger_out
		input  wire [3:0]  pio_1_external_connection_export     //  pio_1_external_connection.export
	);

	wire          altpll_0_c0_clk;                                                                                                // altpll_0:c0 -> [PWM0:csi_I_clk, PWM0_avalon_slave_translator:clk, PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:clk, PWM0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, PWM1:csi_I_clk, PWM1_avalon_slave_translator:clk, PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:clk, PWM1_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, PWM2:csi_I_clk, PWM2_avalon_slave_translator:clk, PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:clk, PWM2_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, PWM3:csi_I_clk, PWM3_avalon_slave_translator:clk, PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:clk, PWM3_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Ultrasound0:clk, Ultrasound0_avalon_slave_0_translator:clk, Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Ultrasound1:clk, Ultrasound1_avalon_slave_0_translator:clk, Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Ultrasound2:clk, Ultrasound2_avalon_slave_0_translator:clk, Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Ultrasound3:clk, Ultrasound3_avalon_slave_0_translator:clk, Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Ultrasound4:clk, Ultrasound4_avalon_slave_0_translator:clk, Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Ultrasound5:clk, Ultrasound5_avalon_slave_0_translator:clk, Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, addr_router:clk, addr_router_001:clk, burst_adapter:clk, cmd_xbar_demux:clk, cmd_xbar_demux_001:clk, cmd_xbar_mux:clk, cmd_xbar_mux_001:clk, cmd_xbar_mux_002:clk, cmd_xbar_mux_003:clk, crosser:in_clk, crosser_001:out_clk, encoder0:clk, encoder0_avalon_slave_0_translator:clk, encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, encoder1:clk, encoder1_avalon_slave_0_translator:clk, encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, epcs_flash_controller_0:clk, epcs_flash_controller_0_epcs_control_port_translator:clk, epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:clk, epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, id_router:clk, id_router_001:clk, id_router_002:clk, id_router_003:clk, id_router_004:clk, id_router_005:clk, id_router_006:clk, id_router_007:clk, id_router_008:clk, id_router_009:clk, id_router_010:clk, id_router_012:clk, id_router_013:clk, id_router_014:clk, id_router_015:clk, id_router_016:clk, id_router_017:clk, id_router_018:clk, id_router_019:clk, id_router_020:clk, id_router_021:clk, id_router_022:clk, id_router_023:clk, id_router_024:clk, id_router_025:clk, irq_mapper:clk, jtag_uart_0:clk, jtag_uart_0_avalon_jtag_slave_translator:clk, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:clk, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, key:clk, key_s1_translator:clk, key_s1_translator_avalon_universal_slave_0_agent:clk, key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, led:clk, led_s1_translator:clk, led_s1_translator_avalon_universal_slave_0_agent:clk, led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, nios2_qsys_0:clk, nios2_qsys_0_data_master_translator:clk, nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:clk, nios2_qsys_0_instruction_master_translator:clk, nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:clk, nios2_qsys_0_jtag_debug_module_translator:clk, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:clk, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, onchip_memory2_0:clk, onchip_memory2_0_s1_translator:clk, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:clk, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, performance_counter:clk, performance_counter_control_slave_translator:clk, performance_counter_control_slave_translator_avalon_universal_slave_0_agent:clk, performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_0:clk, pio_0_s1_translator:clk, pio_0_s1_translator_avalon_universal_slave_0_agent:clk, pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_1:clk, pio_1_s1_translator:clk, pio_1_s1_translator_avalon_universal_slave_0_agent:clk, pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_003:clk, rsp_xbar_demux_004:clk, rsp_xbar_demux_005:clk, rsp_xbar_demux_006:clk, rsp_xbar_demux_007:clk, rsp_xbar_demux_008:clk, rsp_xbar_demux_009:clk, rsp_xbar_demux_010:clk, rsp_xbar_demux_012:clk, rsp_xbar_demux_013:clk, rsp_xbar_demux_014:clk, rsp_xbar_demux_015:clk, rsp_xbar_demux_016:clk, rsp_xbar_demux_017:clk, rsp_xbar_demux_018:clk, rsp_xbar_demux_019:clk, rsp_xbar_demux_020:clk, rsp_xbar_demux_021:clk, rsp_xbar_demux_022:clk, rsp_xbar_demux_023:clk, rsp_xbar_demux_024:clk, rsp_xbar_demux_025:clk, rsp_xbar_mux:clk, rsp_xbar_mux_001:clk, rst_controller:clk, rst_controller_001:clk, sdram:clk, sdram_s1_translator:clk, sdram_s1_translator_avalon_universal_slave_0_agent:clk, sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, sw:clk, sw_s1_translator:clk, sw_s1_translator_avalon_universal_slave_0_agent:clk, sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, timer:clk, timer_s1_translator:clk, timer_s1_translator_avalon_universal_slave_0_agent:clk, timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, uart_0:clk, uart_0_s1_translator:clk, uart_0_s1_translator_avalon_universal_slave_0_agent:clk, uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, width_adapter:clk, width_adapter_001:clk]
	wire          altpll_0_c2_clk;                                                                                                // altpll_0:c2 -> [adc_spi_read:clk, adc_spi_read_slave_translator:clk, adc_spi_read_slave_translator_avalon_universal_slave_0_agent:clk, adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, crosser:out_clk, crosser_001:in_clk, id_router_011:clk, rsp_xbar_demux_011:clk, rst_controller_003:clk]
	wire          nios2_qsys_0_instruction_master_waitrequest;                                                                    // nios2_qsys_0_instruction_master_translator:av_waitrequest -> nios2_qsys_0:i_waitrequest
	wire   [25:0] nios2_qsys_0_instruction_master_address;                                                                        // nios2_qsys_0:i_address -> nios2_qsys_0_instruction_master_translator:av_address
	wire          nios2_qsys_0_instruction_master_read;                                                                           // nios2_qsys_0:i_read -> nios2_qsys_0_instruction_master_translator:av_read
	wire   [31:0] nios2_qsys_0_instruction_master_readdata;                                                                       // nios2_qsys_0_instruction_master_translator:av_readdata -> nios2_qsys_0:i_readdata
	wire          nios2_qsys_0_data_master_waitrequest;                                                                           // nios2_qsys_0_data_master_translator:av_waitrequest -> nios2_qsys_0:d_waitrequest
	wire   [31:0] nios2_qsys_0_data_master_writedata;                                                                             // nios2_qsys_0:d_writedata -> nios2_qsys_0_data_master_translator:av_writedata
	wire   [25:0] nios2_qsys_0_data_master_address;                                                                               // nios2_qsys_0:d_address -> nios2_qsys_0_data_master_translator:av_address
	wire          nios2_qsys_0_data_master_write;                                                                                 // nios2_qsys_0:d_write -> nios2_qsys_0_data_master_translator:av_write
	wire          nios2_qsys_0_data_master_read;                                                                                  // nios2_qsys_0:d_read -> nios2_qsys_0_data_master_translator:av_read
	wire   [31:0] nios2_qsys_0_data_master_readdata;                                                                              // nios2_qsys_0_data_master_translator:av_readdata -> nios2_qsys_0:d_readdata
	wire          nios2_qsys_0_data_master_debugaccess;                                                                           // nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> nios2_qsys_0_data_master_translator:av_debugaccess
	wire    [3:0] nios2_qsys_0_data_master_byteenable;                                                                            // nios2_qsys_0:d_byteenable -> nios2_qsys_0_data_master_translator:av_byteenable
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest;                                      // nios2_qsys_0:jtag_debug_module_waitrequest -> nios2_qsys_0_jtag_debug_module_translator:av_waitrequest
	wire   [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                        // nios2_qsys_0_jtag_debug_module_translator:av_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	wire    [8:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address;                                          // nios2_qsys_0_jtag_debug_module_translator:av_address -> nios2_qsys_0:jtag_debug_module_address
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write;                                            // nios2_qsys_0_jtag_debug_module_translator:av_write -> nios2_qsys_0:jtag_debug_module_write
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_read;                                             // nios2_qsys_0_jtag_debug_module_translator:av_read -> nios2_qsys_0:jtag_debug_module_read
	wire   [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                         // nios2_qsys_0:jtag_debug_module_readdata -> nios2_qsys_0_jtag_debug_module_translator:av_readdata
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                      // nios2_qsys_0_jtag_debug_module_translator:av_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	wire    [3:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                       // nios2_qsys_0_jtag_debug_module_translator:av_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	wire          sdram_s1_translator_avalon_anti_slave_0_waitrequest;                                                            // sdram:za_waitrequest -> sdram_s1_translator:av_waitrequest
	wire   [15:0] sdram_s1_translator_avalon_anti_slave_0_writedata;                                                              // sdram_s1_translator:av_writedata -> sdram:az_data
	wire   [23:0] sdram_s1_translator_avalon_anti_slave_0_address;                                                                // sdram_s1_translator:av_address -> sdram:az_addr
	wire          sdram_s1_translator_avalon_anti_slave_0_chipselect;                                                             // sdram_s1_translator:av_chipselect -> sdram:az_cs
	wire          sdram_s1_translator_avalon_anti_slave_0_write;                                                                  // sdram_s1_translator:av_write -> sdram:az_wr_n
	wire          sdram_s1_translator_avalon_anti_slave_0_read;                                                                   // sdram_s1_translator:av_read -> sdram:az_rd_n
	wire   [15:0] sdram_s1_translator_avalon_anti_slave_0_readdata;                                                               // sdram:za_data -> sdram_s1_translator:av_readdata
	wire          sdram_s1_translator_avalon_anti_slave_0_readdatavalid;                                                          // sdram:za_valid -> sdram_s1_translator:av_readdatavalid
	wire    [1:0] sdram_s1_translator_avalon_anti_slave_0_byteenable;                                                             // sdram_s1_translator:av_byteenable -> sdram:az_be_n
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata;                                                   // onchip_memory2_0_s1_translator:av_writedata -> onchip_memory2_0:writedata
	wire   [11:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_address;                                                     // onchip_memory2_0_s1_translator:av_address -> onchip_memory2_0:address
	wire          onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect;                                                  // onchip_memory2_0_s1_translator:av_chipselect -> onchip_memory2_0:chipselect
	wire          onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken;                                                       // onchip_memory2_0_s1_translator:av_clken -> onchip_memory2_0:clken
	wire          onchip_memory2_0_s1_translator_avalon_anti_slave_0_write;                                                       // onchip_memory2_0_s1_translator:av_write -> onchip_memory2_0:write
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata;                                                    // onchip_memory2_0:readdata -> onchip_memory2_0_s1_translator:av_readdata
	wire    [3:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable;                                                  // onchip_memory2_0_s1_translator:av_byteenable -> onchip_memory2_0:byteenable
	wire   [31:0] epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_writedata;                             // epcs_flash_controller_0_epcs_control_port_translator:av_writedata -> epcs_flash_controller_0:writedata
	wire    [8:0] epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_address;                               // epcs_flash_controller_0_epcs_control_port_translator:av_address -> epcs_flash_controller_0:address
	wire          epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_chipselect;                            // epcs_flash_controller_0_epcs_control_port_translator:av_chipselect -> epcs_flash_controller_0:chipselect
	wire          epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_write;                                 // epcs_flash_controller_0_epcs_control_port_translator:av_write -> epcs_flash_controller_0:write_n
	wire          epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_read;                                  // epcs_flash_controller_0_epcs_control_port_translator:av_read -> epcs_flash_controller_0:read_n
	wire   [31:0] epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_readdata;                              // epcs_flash_controller_0:readdata -> epcs_flash_controller_0_epcs_control_port_translator:av_readdata
	wire   [31:0] led_s1_translator_avalon_anti_slave_0_writedata;                                                                // led_s1_translator:av_writedata -> led:writedata
	wire    [1:0] led_s1_translator_avalon_anti_slave_0_address;                                                                  // led_s1_translator:av_address -> led:address
	wire          led_s1_translator_avalon_anti_slave_0_chipselect;                                                               // led_s1_translator:av_chipselect -> led:chipselect
	wire          led_s1_translator_avalon_anti_slave_0_write;                                                                    // led_s1_translator:av_write -> led:write_n
	wire   [31:0] led_s1_translator_avalon_anti_slave_0_readdata;                                                                 // led:readdata -> led_s1_translator:av_readdata
	wire   [31:0] key_s1_translator_avalon_anti_slave_0_writedata;                                                                // key_s1_translator:av_writedata -> key:writedata
	wire    [1:0] key_s1_translator_avalon_anti_slave_0_address;                                                                  // key_s1_translator:av_address -> key:address
	wire          key_s1_translator_avalon_anti_slave_0_chipselect;                                                               // key_s1_translator:av_chipselect -> key:chipselect
	wire          key_s1_translator_avalon_anti_slave_0_write;                                                                    // key_s1_translator:av_write -> key:write_n
	wire   [31:0] key_s1_translator_avalon_anti_slave_0_readdata;                                                                 // key:readdata -> key_s1_translator:av_readdata
	wire   [31:0] sw_s1_translator_avalon_anti_slave_0_writedata;                                                                 // sw_s1_translator:av_writedata -> sw:writedata
	wire    [1:0] sw_s1_translator_avalon_anti_slave_0_address;                                                                   // sw_s1_translator:av_address -> sw:address
	wire          sw_s1_translator_avalon_anti_slave_0_chipselect;                                                                // sw_s1_translator:av_chipselect -> sw:chipselect
	wire          sw_s1_translator_avalon_anti_slave_0_write;                                                                     // sw_s1_translator:av_write -> sw:write_n
	wire   [31:0] sw_s1_translator_avalon_anti_slave_0_readdata;                                                                  // sw:readdata -> sw_s1_translator:av_readdata
	wire   [15:0] timer_s1_translator_avalon_anti_slave_0_writedata;                                                              // timer_s1_translator:av_writedata -> timer:writedata
	wire    [2:0] timer_s1_translator_avalon_anti_slave_0_address;                                                                // timer_s1_translator:av_address -> timer:address
	wire          timer_s1_translator_avalon_anti_slave_0_chipselect;                                                             // timer_s1_translator:av_chipselect -> timer:chipselect
	wire          timer_s1_translator_avalon_anti_slave_0_write;                                                                  // timer_s1_translator:av_write -> timer:write_n
	wire   [15:0] timer_s1_translator_avalon_anti_slave_0_readdata;                                                               // timer:readdata -> timer_s1_translator:av_readdata
	wire   [31:0] performance_counter_control_slave_translator_avalon_anti_slave_0_writedata;                                     // performance_counter_control_slave_translator:av_writedata -> performance_counter:writedata
	wire    [3:0] performance_counter_control_slave_translator_avalon_anti_slave_0_address;                                       // performance_counter_control_slave_translator:av_address -> performance_counter:address
	wire          performance_counter_control_slave_translator_avalon_anti_slave_0_write;                                         // performance_counter_control_slave_translator:av_write -> performance_counter:write
	wire   [31:0] performance_counter_control_slave_translator_avalon_anti_slave_0_readdata;                                      // performance_counter:readdata -> performance_counter_control_slave_translator:av_readdata
	wire          performance_counter_control_slave_translator_avalon_anti_slave_0_begintransfer;                                 // performance_counter_control_slave_translator:av_begintransfer -> performance_counter:begintransfer
	wire   [31:0] ultrasound0_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                            // Ultrasound0_avalon_slave_0_translator:av_writedata -> Ultrasound0:writedata
	wire    [1:0] ultrasound0_avalon_slave_0_translator_avalon_anti_slave_0_address;                                              // Ultrasound0_avalon_slave_0_translator:av_address -> Ultrasound0:address
	wire          ultrasound0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                                           // Ultrasound0_avalon_slave_0_translator:av_chipselect -> Ultrasound0:chipselect
	wire          ultrasound0_avalon_slave_0_translator_avalon_anti_slave_0_write;                                                // Ultrasound0_avalon_slave_0_translator:av_write -> Ultrasound0:write
	wire          ultrasound0_avalon_slave_0_translator_avalon_anti_slave_0_read;                                                 // Ultrasound0_avalon_slave_0_translator:av_read -> Ultrasound0:read
	wire   [31:0] ultrasound0_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                             // Ultrasound0:readdata -> Ultrasound0_avalon_slave_0_translator:av_readdata
	wire    [3:0] ultrasound0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable;                                           // Ultrasound0_avalon_slave_0_translator:av_byteenable -> Ultrasound0:byteenable
	wire   [31:0] ultrasound1_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                            // Ultrasound1_avalon_slave_0_translator:av_writedata -> Ultrasound1:writedata
	wire    [1:0] ultrasound1_avalon_slave_0_translator_avalon_anti_slave_0_address;                                              // Ultrasound1_avalon_slave_0_translator:av_address -> Ultrasound1:address
	wire          ultrasound1_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                                           // Ultrasound1_avalon_slave_0_translator:av_chipselect -> Ultrasound1:chipselect
	wire          ultrasound1_avalon_slave_0_translator_avalon_anti_slave_0_write;                                                // Ultrasound1_avalon_slave_0_translator:av_write -> Ultrasound1:write
	wire          ultrasound1_avalon_slave_0_translator_avalon_anti_slave_0_read;                                                 // Ultrasound1_avalon_slave_0_translator:av_read -> Ultrasound1:read
	wire   [31:0] ultrasound1_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                             // Ultrasound1:readdata -> Ultrasound1_avalon_slave_0_translator:av_readdata
	wire    [3:0] ultrasound1_avalon_slave_0_translator_avalon_anti_slave_0_byteenable;                                           // Ultrasound1_avalon_slave_0_translator:av_byteenable -> Ultrasound1:byteenable
	wire   [15:0] adc_spi_read_slave_translator_avalon_anti_slave_0_writedata;                                                    // adc_spi_read_slave_translator:av_writedata -> adc_spi_read:s_writedata
	wire          adc_spi_read_slave_translator_avalon_anti_slave_0_chipselect;                                                   // adc_spi_read_slave_translator:av_chipselect -> adc_spi_read:s_chipselect
	wire          adc_spi_read_slave_translator_avalon_anti_slave_0_write;                                                        // adc_spi_read_slave_translator:av_write -> adc_spi_read:s_write
	wire          adc_spi_read_slave_translator_avalon_anti_slave_0_read;                                                         // adc_spi_read_slave_translator:av_read -> adc_spi_read:s_read
	wire   [15:0] adc_spi_read_slave_translator_avalon_anti_slave_0_readdata;                                                     // adc_spi_read:s_readdata -> adc_spi_read_slave_translator:av_readdata
	wire   [31:0] pwm0_avalon_slave_translator_avalon_anti_slave_0_writedata;                                                     // PWM0_avalon_slave_translator:av_writedata -> PWM0:avs_I_wr_data
	wire    [2:0] pwm0_avalon_slave_translator_avalon_anti_slave_0_address;                                                       // PWM0_avalon_slave_translator:av_address -> PWM0:avs_address
	wire          pwm0_avalon_slave_translator_avalon_anti_slave_0_chipselect;                                                    // PWM0_avalon_slave_translator:av_chipselect -> PWM0:avs_I_cs
	wire          pwm0_avalon_slave_translator_avalon_anti_slave_0_write;                                                         // PWM0_avalon_slave_translator:av_write -> PWM0:avs_write
	wire   [31:0] pwm1_avalon_slave_translator_avalon_anti_slave_0_writedata;                                                     // PWM1_avalon_slave_translator:av_writedata -> PWM1:avs_I_wr_data
	wire    [2:0] pwm1_avalon_slave_translator_avalon_anti_slave_0_address;                                                       // PWM1_avalon_slave_translator:av_address -> PWM1:avs_address
	wire          pwm1_avalon_slave_translator_avalon_anti_slave_0_chipselect;                                                    // PWM1_avalon_slave_translator:av_chipselect -> PWM1:avs_I_cs
	wire          pwm1_avalon_slave_translator_avalon_anti_slave_0_write;                                                         // PWM1_avalon_slave_translator:av_write -> PWM1:avs_write
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                                       // jtag_uart_0:av_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                                         // jtag_uart_0_avalon_jtag_slave_translator:av_writedata -> jtag_uart_0:av_writedata
	wire    [0:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                           // jtag_uart_0_avalon_jtag_slave_translator:av_address -> jtag_uart_0:av_address
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                                        // jtag_uart_0_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_0:av_chipselect
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                             // jtag_uart_0_avalon_jtag_slave_translator:av_write -> jtag_uart_0:av_write_n
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                              // jtag_uart_0_avalon_jtag_slave_translator:av_read -> jtag_uart_0:av_read_n
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                                          // jtag_uart_0:av_readdata -> jtag_uart_0_avalon_jtag_slave_translator:av_readdata
	wire   [31:0] encoder0_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                               // encoder0_avalon_slave_0_translator:av_writedata -> encoder0:writedata
	wire    [1:0] encoder0_avalon_slave_0_translator_avalon_anti_slave_0_address;                                                 // encoder0_avalon_slave_0_translator:av_address -> encoder0:address
	wire          encoder0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                                              // encoder0_avalon_slave_0_translator:av_chipselect -> encoder0:chipselect
	wire          encoder0_avalon_slave_0_translator_avalon_anti_slave_0_write;                                                   // encoder0_avalon_slave_0_translator:av_write -> encoder0:write
	wire          encoder0_avalon_slave_0_translator_avalon_anti_slave_0_read;                                                    // encoder0_avalon_slave_0_translator:av_read -> encoder0:read
	wire   [31:0] encoder0_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                                // encoder0:readdata -> encoder0_avalon_slave_0_translator:av_readdata
	wire    [3:0] encoder0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable;                                              // encoder0_avalon_slave_0_translator:av_byteenable -> encoder0:byteenable
	wire   [31:0] encoder1_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                               // encoder1_avalon_slave_0_translator:av_writedata -> encoder1:writedata
	wire    [1:0] encoder1_avalon_slave_0_translator_avalon_anti_slave_0_address;                                                 // encoder1_avalon_slave_0_translator:av_address -> encoder1:address
	wire          encoder1_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                                              // encoder1_avalon_slave_0_translator:av_chipselect -> encoder1:chipselect
	wire          encoder1_avalon_slave_0_translator_avalon_anti_slave_0_write;                                                   // encoder1_avalon_slave_0_translator:av_write -> encoder1:write
	wire          encoder1_avalon_slave_0_translator_avalon_anti_slave_0_read;                                                    // encoder1_avalon_slave_0_translator:av_read -> encoder1:read
	wire   [31:0] encoder1_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                                // encoder1:readdata -> encoder1_avalon_slave_0_translator:av_readdata
	wire    [3:0] encoder1_avalon_slave_0_translator_avalon_anti_slave_0_byteenable;                                              // encoder1_avalon_slave_0_translator:av_byteenable -> encoder1:byteenable
	wire   [31:0] pio_0_s1_translator_avalon_anti_slave_0_writedata;                                                              // pio_0_s1_translator:av_writedata -> pio_0:writedata
	wire    [1:0] pio_0_s1_translator_avalon_anti_slave_0_address;                                                                // pio_0_s1_translator:av_address -> pio_0:address
	wire          pio_0_s1_translator_avalon_anti_slave_0_chipselect;                                                             // pio_0_s1_translator:av_chipselect -> pio_0:chipselect
	wire          pio_0_s1_translator_avalon_anti_slave_0_write;                                                                  // pio_0_s1_translator:av_write -> pio_0:write_n
	wire   [31:0] pio_0_s1_translator_avalon_anti_slave_0_readdata;                                                               // pio_0:readdata -> pio_0_s1_translator:av_readdata
	wire   [15:0] uart_0_s1_translator_avalon_anti_slave_0_writedata;                                                             // uart_0_s1_translator:av_writedata -> uart_0:writedata
	wire    [2:0] uart_0_s1_translator_avalon_anti_slave_0_address;                                                               // uart_0_s1_translator:av_address -> uart_0:address
	wire          uart_0_s1_translator_avalon_anti_slave_0_chipselect;                                                            // uart_0_s1_translator:av_chipselect -> uart_0:chipselect
	wire          uart_0_s1_translator_avalon_anti_slave_0_write;                                                                 // uart_0_s1_translator:av_write -> uart_0:write_n
	wire          uart_0_s1_translator_avalon_anti_slave_0_read;                                                                  // uart_0_s1_translator:av_read -> uart_0:read_n
	wire   [15:0] uart_0_s1_translator_avalon_anti_slave_0_readdata;                                                              // uart_0:readdata -> uart_0_s1_translator:av_readdata
	wire          uart_0_s1_translator_avalon_anti_slave_0_begintransfer;                                                         // uart_0_s1_translator:av_begintransfer -> uart_0:begintransfer
	wire   [31:0] ultrasound2_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                            // Ultrasound2_avalon_slave_0_translator:av_writedata -> Ultrasound2:writedata
	wire    [1:0] ultrasound2_avalon_slave_0_translator_avalon_anti_slave_0_address;                                              // Ultrasound2_avalon_slave_0_translator:av_address -> Ultrasound2:address
	wire          ultrasound2_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                                           // Ultrasound2_avalon_slave_0_translator:av_chipselect -> Ultrasound2:chipselect
	wire          ultrasound2_avalon_slave_0_translator_avalon_anti_slave_0_write;                                                // Ultrasound2_avalon_slave_0_translator:av_write -> Ultrasound2:write
	wire          ultrasound2_avalon_slave_0_translator_avalon_anti_slave_0_read;                                                 // Ultrasound2_avalon_slave_0_translator:av_read -> Ultrasound2:read
	wire   [31:0] ultrasound2_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                             // Ultrasound2:readdata -> Ultrasound2_avalon_slave_0_translator:av_readdata
	wire    [3:0] ultrasound2_avalon_slave_0_translator_avalon_anti_slave_0_byteenable;                                           // Ultrasound2_avalon_slave_0_translator:av_byteenable -> Ultrasound2:byteenable
	wire   [31:0] ultrasound3_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                            // Ultrasound3_avalon_slave_0_translator:av_writedata -> Ultrasound3:writedata
	wire    [1:0] ultrasound3_avalon_slave_0_translator_avalon_anti_slave_0_address;                                              // Ultrasound3_avalon_slave_0_translator:av_address -> Ultrasound3:address
	wire          ultrasound3_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                                           // Ultrasound3_avalon_slave_0_translator:av_chipselect -> Ultrasound3:chipselect
	wire          ultrasound3_avalon_slave_0_translator_avalon_anti_slave_0_write;                                                // Ultrasound3_avalon_slave_0_translator:av_write -> Ultrasound3:write
	wire          ultrasound3_avalon_slave_0_translator_avalon_anti_slave_0_read;                                                 // Ultrasound3_avalon_slave_0_translator:av_read -> Ultrasound3:read
	wire   [31:0] ultrasound3_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                             // Ultrasound3:readdata -> Ultrasound3_avalon_slave_0_translator:av_readdata
	wire    [3:0] ultrasound3_avalon_slave_0_translator_avalon_anti_slave_0_byteenable;                                           // Ultrasound3_avalon_slave_0_translator:av_byteenable -> Ultrasound3:byteenable
	wire   [31:0] ultrasound4_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                            // Ultrasound4_avalon_slave_0_translator:av_writedata -> Ultrasound4:writedata
	wire    [1:0] ultrasound4_avalon_slave_0_translator_avalon_anti_slave_0_address;                                              // Ultrasound4_avalon_slave_0_translator:av_address -> Ultrasound4:address
	wire          ultrasound4_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                                           // Ultrasound4_avalon_slave_0_translator:av_chipselect -> Ultrasound4:chipselect
	wire          ultrasound4_avalon_slave_0_translator_avalon_anti_slave_0_write;                                                // Ultrasound4_avalon_slave_0_translator:av_write -> Ultrasound4:write
	wire          ultrasound4_avalon_slave_0_translator_avalon_anti_slave_0_read;                                                 // Ultrasound4_avalon_slave_0_translator:av_read -> Ultrasound4:read
	wire   [31:0] ultrasound4_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                             // Ultrasound4:readdata -> Ultrasound4_avalon_slave_0_translator:av_readdata
	wire    [3:0] ultrasound4_avalon_slave_0_translator_avalon_anti_slave_0_byteenable;                                           // Ultrasound4_avalon_slave_0_translator:av_byteenable -> Ultrasound4:byteenable
	wire   [31:0] ultrasound5_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                            // Ultrasound5_avalon_slave_0_translator:av_writedata -> Ultrasound5:writedata
	wire    [1:0] ultrasound5_avalon_slave_0_translator_avalon_anti_slave_0_address;                                              // Ultrasound5_avalon_slave_0_translator:av_address -> Ultrasound5:address
	wire          ultrasound5_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                                           // Ultrasound5_avalon_slave_0_translator:av_chipselect -> Ultrasound5:chipselect
	wire          ultrasound5_avalon_slave_0_translator_avalon_anti_slave_0_write;                                                // Ultrasound5_avalon_slave_0_translator:av_write -> Ultrasound5:write
	wire          ultrasound5_avalon_slave_0_translator_avalon_anti_slave_0_read;                                                 // Ultrasound5_avalon_slave_0_translator:av_read -> Ultrasound5:read
	wire   [31:0] ultrasound5_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                             // Ultrasound5:readdata -> Ultrasound5_avalon_slave_0_translator:av_readdata
	wire    [3:0] ultrasound5_avalon_slave_0_translator_avalon_anti_slave_0_byteenable;                                           // Ultrasound5_avalon_slave_0_translator:av_byteenable -> Ultrasound5:byteenable
	wire   [31:0] pwm2_avalon_slave_translator_avalon_anti_slave_0_writedata;                                                     // PWM2_avalon_slave_translator:av_writedata -> PWM2:avs_I_wr_data
	wire    [2:0] pwm2_avalon_slave_translator_avalon_anti_slave_0_address;                                                       // PWM2_avalon_slave_translator:av_address -> PWM2:avs_address
	wire          pwm2_avalon_slave_translator_avalon_anti_slave_0_chipselect;                                                    // PWM2_avalon_slave_translator:av_chipselect -> PWM2:avs_I_cs
	wire          pwm2_avalon_slave_translator_avalon_anti_slave_0_write;                                                         // PWM2_avalon_slave_translator:av_write -> PWM2:avs_write
	wire   [31:0] pwm3_avalon_slave_translator_avalon_anti_slave_0_writedata;                                                     // PWM3_avalon_slave_translator:av_writedata -> PWM3:avs_I_wr_data
	wire    [2:0] pwm3_avalon_slave_translator_avalon_anti_slave_0_address;                                                       // PWM3_avalon_slave_translator:av_address -> PWM3:avs_address
	wire          pwm3_avalon_slave_translator_avalon_anti_slave_0_chipselect;                                                    // PWM3_avalon_slave_translator:av_chipselect -> PWM3:avs_I_cs
	wire          pwm3_avalon_slave_translator_avalon_anti_slave_0_write;                                                         // PWM3_avalon_slave_translator:av_write -> PWM3:avs_write
	wire    [1:0] pio_1_s1_translator_avalon_anti_slave_0_address;                                                                // pio_1_s1_translator:av_address -> pio_1:address
	wire   [31:0] pio_1_s1_translator_avalon_anti_slave_0_readdata;                                                               // pio_1:readdata -> pio_1_s1_translator:av_readdata
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest;                               // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_0_instruction_master_translator:uav_waitrequest
	wire    [2:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount;                                // nios2_qsys_0_instruction_master_translator:uav_burstcount -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata;                                 // nios2_qsys_0_instruction_master_translator:uav_writedata -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [25:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address;                                   // nios2_qsys_0_instruction_master_translator:uav_address -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock;                                      // nios2_qsys_0_instruction_master_translator:uav_lock -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write;                                     // nios2_qsys_0_instruction_master_translator:uav_write -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read;                                      // nios2_qsys_0_instruction_master_translator:uav_read -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata;                                  // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_0_instruction_master_translator:uav_readdata
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess;                               // nios2_qsys_0_instruction_master_translator:uav_debugaccess -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable;                                // nios2_qsys_0_instruction_master_translator:uav_byteenable -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid;                             // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_0_instruction_master_translator:uav_readdatavalid
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest;                                      // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_0_data_master_translator:uav_waitrequest
	wire    [2:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount;                                       // nios2_qsys_0_data_master_translator:uav_burstcount -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata;                                        // nios2_qsys_0_data_master_translator:uav_writedata -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [25:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_address;                                          // nios2_qsys_0_data_master_translator:uav_address -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock;                                             // nios2_qsys_0_data_master_translator:uav_lock -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_write;                                            // nios2_qsys_0_data_master_translator:uav_write -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_read;                                             // nios2_qsys_0_data_master_translator:uav_read -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata;                                         // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_0_data_master_translator:uav_readdata
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess;                                      // nios2_qsys_0_data_master_translator:uav_debugaccess -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable;                                       // nios2_qsys_0_data_master_translator:uav_byteenable -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid;                                    // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_0_data_master_translator:uav_readdatavalid
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // nios2_qsys_0_jtag_debug_module_translator:uav_waitrequest -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2_qsys_0_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                          // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2_qsys_0_jtag_debug_module_translator:uav_writedata
	wire   [25:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                            // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2_qsys_0_jtag_debug_module_translator:uav_address
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                              // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2_qsys_0_jtag_debug_module_translator:uav_write
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                               // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2_qsys_0_jtag_debug_module_translator:uav_lock
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                               // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2_qsys_0_jtag_debug_module_translator:uav_read
	wire   [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                           // nios2_qsys_0_jtag_debug_module_translator:uav_readdata -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // nios2_qsys_0_jtag_debug_module_translator:uav_readdatavalid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2_qsys_0_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2_qsys_0_jtag_debug_module_translator:uav_byteenable
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                        // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                              // sdram_s1_translator:uav_waitrequest -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                               // sdram_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_s1_translator:uav_burstcount
	wire   [15:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                // sdram_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_s1_translator:uav_writedata
	wire   [25:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                  // sdram_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdram_s1_translator:uav_address
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                    // sdram_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdram_s1_translator:uav_write
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                     // sdram_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_s1_translator:uav_lock
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                     // sdram_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdram_s1_translator:uav_read
	wire   [15:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                 // sdram_s1_translator:uav_readdata -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                            // sdram_s1_translator:uav_readdatavalid -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                              // sdram_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_s1_translator:uav_debugaccess
	wire    [1:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                               // sdram_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_s1_translator:uav_byteenable
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                       // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                             // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                     // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [85:0] sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                              // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                             // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                    // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                          // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                  // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [85:0] sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                           // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                          // sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                        // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [17:0] sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                         // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                        // sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                                        // sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [17:0] sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                         // sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                                        // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // onchip_memory2_0_s1_translator:uav_waitrequest -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> onchip_memory2_0_s1_translator:uav_burstcount
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> onchip_memory2_0_s1_translator:uav_writedata
	wire   [25:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                       // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> onchip_memory2_0_s1_translator:uav_address
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                         // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> onchip_memory2_0_s1_translator:uav_write
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                          // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> onchip_memory2_0_s1_translator:uav_lock
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                          // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> onchip_memory2_0_s1_translator:uav_read
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // onchip_memory2_0_s1_translator:uav_readdata -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // onchip_memory2_0_s1_translator:uav_readdatavalid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> onchip_memory2_0_s1_translator:uav_debugaccess
	wire    [3:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> onchip_memory2_0_s1_translator:uav_byteenable
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // epcs_flash_controller_0_epcs_control_port_translator:uav_waitrequest -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount;              // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_burstcount -> epcs_flash_controller_0_epcs_control_port_translator:uav_burstcount
	wire   [31:0] epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_writedata;               // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_writedata -> epcs_flash_controller_0_epcs_control_port_translator:uav_writedata
	wire   [25:0] epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_address;                 // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_address -> epcs_flash_controller_0_epcs_control_port_translator:uav_address
	wire          epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_write;                   // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_write -> epcs_flash_controller_0_epcs_control_port_translator:uav_write
	wire          epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_lock;                    // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_lock -> epcs_flash_controller_0_epcs_control_port_translator:uav_lock
	wire          epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_read;                    // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_read -> epcs_flash_controller_0_epcs_control_port_translator:uav_read
	wire   [31:0] epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdata;                // epcs_flash_controller_0_epcs_control_port_translator:uav_readdata -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // epcs_flash_controller_0_epcs_control_port_translator:uav_readdatavalid -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_debugaccess -> epcs_flash_controller_0_epcs_control_port_translator:uav_debugaccess
	wire    [3:0] epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable;              // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_byteenable -> epcs_flash_controller_0_epcs_control_port_translator:uav_byteenable
	wire          epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid;            // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_valid -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_data;             // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_data -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready;            // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_ready -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                // led_s1_translator:uav_waitrequest -> led_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                 // led_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> led_s1_translator:uav_burstcount
	wire   [31:0] led_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                  // led_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> led_s1_translator:uav_writedata
	wire   [25:0] led_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                    // led_s1_translator_avalon_universal_slave_0_agent:m0_address -> led_s1_translator:uav_address
	wire          led_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                      // led_s1_translator_avalon_universal_slave_0_agent:m0_write -> led_s1_translator:uav_write
	wire          led_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                       // led_s1_translator_avalon_universal_slave_0_agent:m0_lock -> led_s1_translator:uav_lock
	wire          led_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                       // led_s1_translator_avalon_universal_slave_0_agent:m0_read -> led_s1_translator:uav_read
	wire   [31:0] led_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                   // led_s1_translator:uav_readdata -> led_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                              // led_s1_translator:uav_readdatavalid -> led_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                // led_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> led_s1_translator:uav_debugaccess
	wire    [3:0] led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                 // led_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> led_s1_translator:uav_byteenable
	wire          led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                         // led_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                               // led_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                       // led_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] led_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                // led_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                               // led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> led_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                      // led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                            // led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                    // led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                             // led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                            // led_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                          // led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                           // led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                          // led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          key_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                // key_s1_translator:uav_waitrequest -> key_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] key_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                 // key_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> key_s1_translator:uav_burstcount
	wire   [31:0] key_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                  // key_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> key_s1_translator:uav_writedata
	wire   [25:0] key_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                    // key_s1_translator_avalon_universal_slave_0_agent:m0_address -> key_s1_translator:uav_address
	wire          key_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                      // key_s1_translator_avalon_universal_slave_0_agent:m0_write -> key_s1_translator:uav_write
	wire          key_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                       // key_s1_translator_avalon_universal_slave_0_agent:m0_lock -> key_s1_translator:uav_lock
	wire          key_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                       // key_s1_translator_avalon_universal_slave_0_agent:m0_read -> key_s1_translator:uav_read
	wire   [31:0] key_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                   // key_s1_translator:uav_readdata -> key_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          key_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                              // key_s1_translator:uav_readdatavalid -> key_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          key_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                // key_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> key_s1_translator:uav_debugaccess
	wire    [3:0] key_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                 // key_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> key_s1_translator:uav_byteenable
	wire          key_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                         // key_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          key_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                               // key_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          key_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                       // key_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] key_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                // key_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          key_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                               // key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> key_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                      // key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> key_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                            // key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> key_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                    // key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> key_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                             // key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> key_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                            // key_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                          // key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                           // key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                          // key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                 // sw_s1_translator:uav_waitrequest -> sw_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                  // sw_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sw_s1_translator:uav_burstcount
	wire   [31:0] sw_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                   // sw_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sw_s1_translator:uav_writedata
	wire   [25:0] sw_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                     // sw_s1_translator_avalon_universal_slave_0_agent:m0_address -> sw_s1_translator:uav_address
	wire          sw_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                       // sw_s1_translator_avalon_universal_slave_0_agent:m0_write -> sw_s1_translator:uav_write
	wire          sw_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                        // sw_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sw_s1_translator:uav_lock
	wire          sw_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                        // sw_s1_translator_avalon_universal_slave_0_agent:m0_read -> sw_s1_translator:uav_read
	wire   [31:0] sw_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                    // sw_s1_translator:uav_readdata -> sw_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                               // sw_s1_translator:uav_readdatavalid -> sw_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                 // sw_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sw_s1_translator:uav_debugaccess
	wire    [3:0] sw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                  // sw_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sw_s1_translator:uav_byteenable
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                          // sw_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                // sw_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                        // sw_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] sw_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                 // sw_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                // sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sw_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                       // sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sw_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                             // sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sw_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                     // sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sw_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                              // sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sw_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                             // sw_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                           // sw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                            // sw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                           // sw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                              // timer_s1_translator:uav_waitrequest -> timer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                               // timer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_s1_translator:uav_burstcount
	wire   [31:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                // timer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_s1_translator:uav_writedata
	wire   [25:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                  // timer_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_s1_translator:uav_address
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                    // timer_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_s1_translator:uav_write
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                     // timer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_s1_translator:uav_lock
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                     // timer_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_s1_translator:uav_read
	wire   [31:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                 // timer_s1_translator:uav_readdata -> timer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                            // timer_s1_translator:uav_readdatavalid -> timer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                              // timer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_s1_translator:uav_debugaccess
	wire    [3:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                               // timer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_s1_translator:uav_byteenable
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                       // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                             // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                     // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                              // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                             // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                    // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                          // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                  // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                           // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                          // timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                        // timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                         // timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                        // timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // performance_counter_control_slave_translator:uav_waitrequest -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> performance_counter_control_slave_translator:uav_burstcount
	wire   [31:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                       // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> performance_counter_control_slave_translator:uav_writedata
	wire   [25:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                         // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> performance_counter_control_slave_translator:uav_address
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                           // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> performance_counter_control_slave_translator:uav_write
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                            // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> performance_counter_control_slave_translator:uav_lock
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                            // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> performance_counter_control_slave_translator:uav_read
	wire   [31:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                        // performance_counter_control_slave_translator:uav_readdata -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // performance_counter_control_slave_translator:uav_readdatavalid -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> performance_counter_control_slave_translator:uav_debugaccess
	wire    [3:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> performance_counter_control_slave_translator:uav_byteenable
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                     // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // Ultrasound0_avalon_slave_0_translator:uav_waitrequest -> Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> Ultrasound0_avalon_slave_0_translator:uav_burstcount
	wire   [31:0] ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                              // Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> Ultrasound0_avalon_slave_0_translator:uav_writedata
	wire   [25:0] ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                                // Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> Ultrasound0_avalon_slave_0_translator:uav_address
	wire          ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                                  // Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> Ultrasound0_avalon_slave_0_translator:uav_write
	wire          ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                                   // Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> Ultrasound0_avalon_slave_0_translator:uav_lock
	wire          ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                                   // Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> Ultrasound0_avalon_slave_0_translator:uav_read
	wire   [31:0] ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                               // Ultrasound0_avalon_slave_0_translator:uav_readdata -> Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // Ultrasound0_avalon_slave_0_translator:uav_readdatavalid -> Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Ultrasound0_avalon_slave_0_translator:uav_debugaccess
	wire    [3:0] ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> Ultrasound0_avalon_slave_0_translator:uav_byteenable
	wire          ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                            // Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // Ultrasound1_avalon_slave_0_translator:uav_waitrequest -> Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> Ultrasound1_avalon_slave_0_translator:uav_burstcount
	wire   [31:0] ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                              // Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> Ultrasound1_avalon_slave_0_translator:uav_writedata
	wire   [25:0] ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                                // Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> Ultrasound1_avalon_slave_0_translator:uav_address
	wire          ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                                  // Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> Ultrasound1_avalon_slave_0_translator:uav_write
	wire          ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                                   // Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> Ultrasound1_avalon_slave_0_translator:uav_lock
	wire          ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                                   // Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> Ultrasound1_avalon_slave_0_translator:uav_read
	wire   [31:0] ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                               // Ultrasound1_avalon_slave_0_translator:uav_readdata -> Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // Ultrasound1_avalon_slave_0_translator:uav_readdatavalid -> Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Ultrasound1_avalon_slave_0_translator:uav_debugaccess
	wire    [3:0] ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> Ultrasound1_avalon_slave_0_translator:uav_byteenable
	wire          ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                            // Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          adc_spi_read_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // adc_spi_read_slave_translator:uav_waitrequest -> adc_spi_read_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] adc_spi_read_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // adc_spi_read_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> adc_spi_read_slave_translator:uav_burstcount
	wire   [31:0] adc_spi_read_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // adc_spi_read_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> adc_spi_read_slave_translator:uav_writedata
	wire   [25:0] adc_spi_read_slave_translator_avalon_universal_slave_0_agent_m0_address;                                        // adc_spi_read_slave_translator_avalon_universal_slave_0_agent:m0_address -> adc_spi_read_slave_translator:uav_address
	wire          adc_spi_read_slave_translator_avalon_universal_slave_0_agent_m0_write;                                          // adc_spi_read_slave_translator_avalon_universal_slave_0_agent:m0_write -> adc_spi_read_slave_translator:uav_write
	wire          adc_spi_read_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                           // adc_spi_read_slave_translator_avalon_universal_slave_0_agent:m0_lock -> adc_spi_read_slave_translator:uav_lock
	wire          adc_spi_read_slave_translator_avalon_universal_slave_0_agent_m0_read;                                           // adc_spi_read_slave_translator_avalon_universal_slave_0_agent:m0_read -> adc_spi_read_slave_translator:uav_read
	wire   [31:0] adc_spi_read_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // adc_spi_read_slave_translator:uav_readdata -> adc_spi_read_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          adc_spi_read_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // adc_spi_read_slave_translator:uav_readdatavalid -> adc_spi_read_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          adc_spi_read_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // adc_spi_read_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> adc_spi_read_slave_translator:uav_debugaccess
	wire    [3:0] adc_spi_read_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // adc_spi_read_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> adc_spi_read_slave_translator:uav_byteenable
	wire          adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // adc_spi_read_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // adc_spi_read_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // adc_spi_read_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // adc_spi_read_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> adc_spi_read_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> adc_spi_read_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> adc_spi_read_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> adc_spi_read_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> adc_spi_read_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // adc_spi_read_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // adc_spi_read_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // adc_spi_read_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> adc_spi_read_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                              // adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> adc_spi_read_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                               // adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> adc_spi_read_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                              // adc_spi_read_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                     // PWM0_avalon_slave_translator:uav_waitrequest -> PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                      // PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> PWM0_avalon_slave_translator:uav_burstcount
	wire   [31:0] pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                       // PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> PWM0_avalon_slave_translator:uav_writedata
	wire   [25:0] pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address;                                         // PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_address -> PWM0_avalon_slave_translator:uav_address
	wire          pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write;                                           // PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_write -> PWM0_avalon_slave_translator:uav_write
	wire          pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                            // PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_lock -> PWM0_avalon_slave_translator:uav_lock
	wire          pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read;                                            // PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_read -> PWM0_avalon_slave_translator:uav_read
	wire   [31:0] pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                        // PWM0_avalon_slave_translator:uav_readdata -> PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                   // PWM0_avalon_slave_translator:uav_readdatavalid -> PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                     // PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> PWM0_avalon_slave_translator:uav_debugaccess
	wire    [3:0] pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                      // PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> PWM0_avalon_slave_translator:uav_byteenable
	wire          pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                              // PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> PWM0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                    // PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> PWM0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                            // PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> PWM0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                     // PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> PWM0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                    // PWM0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                           // PWM0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                 // PWM0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                         // PWM0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                  // PWM0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                 // PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> PWM0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                               // PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                // PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                               // PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                     // PWM1_avalon_slave_translator:uav_waitrequest -> PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                      // PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> PWM1_avalon_slave_translator:uav_burstcount
	wire   [31:0] pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                       // PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> PWM1_avalon_slave_translator:uav_writedata
	wire   [25:0] pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address;                                         // PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:m0_address -> PWM1_avalon_slave_translator:uav_address
	wire          pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write;                                           // PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:m0_write -> PWM1_avalon_slave_translator:uav_write
	wire          pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                            // PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:m0_lock -> PWM1_avalon_slave_translator:uav_lock
	wire          pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read;                                            // PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:m0_read -> PWM1_avalon_slave_translator:uav_read
	wire   [31:0] pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                        // PWM1_avalon_slave_translator:uav_readdata -> PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                   // PWM1_avalon_slave_translator:uav_readdatavalid -> PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                     // PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> PWM1_avalon_slave_translator:uav_debugaccess
	wire    [3:0] pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                      // PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> PWM1_avalon_slave_translator:uav_byteenable
	wire          pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                              // PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> PWM1_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                    // PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> PWM1_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                            // PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> PWM1_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                     // PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> PWM1_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                    // PWM1_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                           // PWM1_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                 // PWM1_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                         // PWM1_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                  // PWM1_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                 // PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> PWM1_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                               // PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                // PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                               // PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                         // jtag_uart_0_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_0_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                           // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_0_avalon_jtag_slave_translator:uav_writedata
	wire   [25:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_0_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_0_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_0_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                                // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_0_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                            // jtag_uart_0_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                       // jtag_uart_0_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_0_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_0_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                  // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                      // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // encoder0_avalon_slave_0_translator:uav_waitrequest -> encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> encoder0_avalon_slave_0_translator:uav_burstcount
	wire   [31:0] encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> encoder0_avalon_slave_0_translator:uav_writedata
	wire   [25:0] encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                                   // encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> encoder0_avalon_slave_0_translator:uav_address
	wire          encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                                     // encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> encoder0_avalon_slave_0_translator:uav_write
	wire          encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                                      // encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> encoder0_avalon_slave_0_translator:uav_lock
	wire          encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                                      // encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> encoder0_avalon_slave_0_translator:uav_read
	wire   [31:0] encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // encoder0_avalon_slave_0_translator:uav_readdata -> encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // encoder0_avalon_slave_0_translator:uav_readdatavalid -> encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> encoder0_avalon_slave_0_translator:uav_debugaccess
	wire    [3:0] encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> encoder0_avalon_slave_0_translator:uav_byteenable
	wire          encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                               // encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // encoder1_avalon_slave_0_translator:uav_waitrequest -> encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> encoder1_avalon_slave_0_translator:uav_burstcount
	wire   [31:0] encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> encoder1_avalon_slave_0_translator:uav_writedata
	wire   [25:0] encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                                   // encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> encoder1_avalon_slave_0_translator:uav_address
	wire          encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                                     // encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> encoder1_avalon_slave_0_translator:uav_write
	wire          encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                                      // encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> encoder1_avalon_slave_0_translator:uav_lock
	wire          encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                                      // encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> encoder1_avalon_slave_0_translator:uav_read
	wire   [31:0] encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // encoder1_avalon_slave_0_translator:uav_readdata -> encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // encoder1_avalon_slave_0_translator:uav_readdatavalid -> encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> encoder1_avalon_slave_0_translator:uav_debugaccess
	wire    [3:0] encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> encoder1_avalon_slave_0_translator:uav_byteenable
	wire          encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                               // encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                              // pio_0_s1_translator:uav_waitrequest -> pio_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pio_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                               // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_0_s1_translator:uav_burstcount
	wire   [31:0] pio_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_0_s1_translator:uav_writedata
	wire   [25:0] pio_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                  // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_0_s1_translator:uav_address
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                    // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_0_s1_translator:uav_write
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                     // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_0_s1_translator:uav_lock
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                     // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_0_s1_translator:uav_read
	wire   [31:0] pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                 // pio_0_s1_translator:uav_readdata -> pio_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                            // pio_0_s1_translator:uav_readdatavalid -> pio_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                              // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_0_s1_translator:uav_debugaccess
	wire    [3:0] pio_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                               // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_0_s1_translator:uav_byteenable
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                       // pio_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                             // pio_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                     // pio_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                              // pio_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                             // pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                    // pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                          // pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                  // pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                           // pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                          // pio_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                        // pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                         // pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                        // pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                             // uart_0_s1_translator:uav_waitrequest -> uart_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] uart_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                              // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> uart_0_s1_translator:uav_burstcount
	wire   [31:0] uart_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                               // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> uart_0_s1_translator:uav_writedata
	wire   [25:0] uart_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                 // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> uart_0_s1_translator:uav_address
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                   // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> uart_0_s1_translator:uav_write
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                    // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> uart_0_s1_translator:uav_lock
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                    // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> uart_0_s1_translator:uav_read
	wire   [31:0] uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                // uart_0_s1_translator:uav_readdata -> uart_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                           // uart_0_s1_translator:uav_readdatavalid -> uart_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                             // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> uart_0_s1_translator:uav_debugaccess
	wire    [3:0] uart_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                              // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> uart_0_s1_translator:uav_byteenable
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                      // uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                            // uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                    // uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                             // uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                            // uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                   // uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                         // uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                 // uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                          // uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                         // uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                       // uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                        // uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                       // uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // Ultrasound2_avalon_slave_0_translator:uav_waitrequest -> Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> Ultrasound2_avalon_slave_0_translator:uav_burstcount
	wire   [31:0] ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                              // Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> Ultrasound2_avalon_slave_0_translator:uav_writedata
	wire   [25:0] ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                                // Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> Ultrasound2_avalon_slave_0_translator:uav_address
	wire          ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                                  // Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> Ultrasound2_avalon_slave_0_translator:uav_write
	wire          ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                                   // Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> Ultrasound2_avalon_slave_0_translator:uav_lock
	wire          ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                                   // Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> Ultrasound2_avalon_slave_0_translator:uav_read
	wire   [31:0] ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                               // Ultrasound2_avalon_slave_0_translator:uav_readdata -> Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // Ultrasound2_avalon_slave_0_translator:uav_readdatavalid -> Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Ultrasound2_avalon_slave_0_translator:uav_debugaccess
	wire    [3:0] ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> Ultrasound2_avalon_slave_0_translator:uav_byteenable
	wire          ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                            // Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // Ultrasound3_avalon_slave_0_translator:uav_waitrequest -> Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> Ultrasound3_avalon_slave_0_translator:uav_burstcount
	wire   [31:0] ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                              // Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> Ultrasound3_avalon_slave_0_translator:uav_writedata
	wire   [25:0] ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                                // Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> Ultrasound3_avalon_slave_0_translator:uav_address
	wire          ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                                  // Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> Ultrasound3_avalon_slave_0_translator:uav_write
	wire          ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                                   // Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> Ultrasound3_avalon_slave_0_translator:uav_lock
	wire          ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                                   // Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> Ultrasound3_avalon_slave_0_translator:uav_read
	wire   [31:0] ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                               // Ultrasound3_avalon_slave_0_translator:uav_readdata -> Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // Ultrasound3_avalon_slave_0_translator:uav_readdatavalid -> Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Ultrasound3_avalon_slave_0_translator:uav_debugaccess
	wire    [3:0] ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> Ultrasound3_avalon_slave_0_translator:uav_byteenable
	wire          ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                            // Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // Ultrasound4_avalon_slave_0_translator:uav_waitrequest -> Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> Ultrasound4_avalon_slave_0_translator:uav_burstcount
	wire   [31:0] ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                              // Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> Ultrasound4_avalon_slave_0_translator:uav_writedata
	wire   [25:0] ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                                // Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> Ultrasound4_avalon_slave_0_translator:uav_address
	wire          ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                                  // Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> Ultrasound4_avalon_slave_0_translator:uav_write
	wire          ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                                   // Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> Ultrasound4_avalon_slave_0_translator:uav_lock
	wire          ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                                   // Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> Ultrasound4_avalon_slave_0_translator:uav_read
	wire   [31:0] ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                               // Ultrasound4_avalon_slave_0_translator:uav_readdata -> Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // Ultrasound4_avalon_slave_0_translator:uav_readdatavalid -> Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Ultrasound4_avalon_slave_0_translator:uav_debugaccess
	wire    [3:0] ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> Ultrasound4_avalon_slave_0_translator:uav_byteenable
	wire          ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                            // Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // Ultrasound5_avalon_slave_0_translator:uav_waitrequest -> Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> Ultrasound5_avalon_slave_0_translator:uav_burstcount
	wire   [31:0] ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                              // Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> Ultrasound5_avalon_slave_0_translator:uav_writedata
	wire   [25:0] ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                                // Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> Ultrasound5_avalon_slave_0_translator:uav_address
	wire          ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                                  // Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> Ultrasound5_avalon_slave_0_translator:uav_write
	wire          ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                                   // Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> Ultrasound5_avalon_slave_0_translator:uav_lock
	wire          ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                                   // Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> Ultrasound5_avalon_slave_0_translator:uav_read
	wire   [31:0] ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                               // Ultrasound5_avalon_slave_0_translator:uav_readdata -> Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // Ultrasound5_avalon_slave_0_translator:uav_readdatavalid -> Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Ultrasound5_avalon_slave_0_translator:uav_debugaccess
	wire    [3:0] ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> Ultrasound5_avalon_slave_0_translator:uav_byteenable
	wire          ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                            // Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                     // PWM2_avalon_slave_translator:uav_waitrequest -> PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                      // PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> PWM2_avalon_slave_translator:uav_burstcount
	wire   [31:0] pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                       // PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> PWM2_avalon_slave_translator:uav_writedata
	wire   [25:0] pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address;                                         // PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:m0_address -> PWM2_avalon_slave_translator:uav_address
	wire          pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write;                                           // PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:m0_write -> PWM2_avalon_slave_translator:uav_write
	wire          pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                            // PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:m0_lock -> PWM2_avalon_slave_translator:uav_lock
	wire          pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read;                                            // PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:m0_read -> PWM2_avalon_slave_translator:uav_read
	wire   [31:0] pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                        // PWM2_avalon_slave_translator:uav_readdata -> PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                   // PWM2_avalon_slave_translator:uav_readdatavalid -> PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                     // PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> PWM2_avalon_slave_translator:uav_debugaccess
	wire    [3:0] pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                      // PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> PWM2_avalon_slave_translator:uav_byteenable
	wire          pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                              // PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> PWM2_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                    // PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> PWM2_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                            // PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> PWM2_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                     // PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> PWM2_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                    // PWM2_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                           // PWM2_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                 // PWM2_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                         // PWM2_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                  // PWM2_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                 // PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> PWM2_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                               // PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                // PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                               // PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                     // PWM3_avalon_slave_translator:uav_waitrequest -> PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                      // PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> PWM3_avalon_slave_translator:uav_burstcount
	wire   [31:0] pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                       // PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> PWM3_avalon_slave_translator:uav_writedata
	wire   [25:0] pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address;                                         // PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:m0_address -> PWM3_avalon_slave_translator:uav_address
	wire          pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write;                                           // PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:m0_write -> PWM3_avalon_slave_translator:uav_write
	wire          pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                            // PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:m0_lock -> PWM3_avalon_slave_translator:uav_lock
	wire          pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read;                                            // PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:m0_read -> PWM3_avalon_slave_translator:uav_read
	wire   [31:0] pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                        // PWM3_avalon_slave_translator:uav_readdata -> PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                   // PWM3_avalon_slave_translator:uav_readdatavalid -> PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                     // PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> PWM3_avalon_slave_translator:uav_debugaccess
	wire    [3:0] pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                      // PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> PWM3_avalon_slave_translator:uav_byteenable
	wire          pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                              // PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> PWM3_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                    // PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> PWM3_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                            // PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> PWM3_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                     // PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> PWM3_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                    // PWM3_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                           // PWM3_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                 // PWM3_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                         // PWM3_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                  // PWM3_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                 // PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> PWM3_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                               // PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                // PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                               // PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                              // pio_1_s1_translator:uav_waitrequest -> pio_1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pio_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                               // pio_1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_1_s1_translator:uav_burstcount
	wire   [31:0] pio_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                // pio_1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_1_s1_translator:uav_writedata
	wire   [25:0] pio_1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                  // pio_1_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_1_s1_translator:uav_address
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                    // pio_1_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_1_s1_translator:uav_write
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                     // pio_1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_1_s1_translator:uav_lock
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                     // pio_1_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_1_s1_translator:uav_read
	wire   [31:0] pio_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                 // pio_1_s1_translator:uav_readdata -> pio_1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                            // pio_1_s1_translator:uav_readdatavalid -> pio_1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                              // pio_1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_1_s1_translator:uav_debugaccess
	wire    [3:0] pio_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                               // pio_1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_1_s1_translator:uav_byteenable
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                       // pio_1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                             // pio_1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                     // pio_1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                              // pio_1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                             // pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                    // pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                          // pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                  // pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                           // pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                          // pio_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                        // pio_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                         // pio_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                        // pio_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                      // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                            // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                    // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [102:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                             // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                            // addr_router:sink_ready -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                             // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid;                                   // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                           // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [102:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data;                                    // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready;                                   // addr_router_001:sink_ready -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                              // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [102:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                               // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router:sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                              // sdram_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                    // sdram_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                            // sdram_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire   [84:0] sdram_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                     // sdram_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                    // id_router_001:sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                         // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [102:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                          // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router_002:sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_valid;                   // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [102:0] epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_data;                    // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_003:sink_ready -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_ready
	wire          led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                // led_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          led_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                      // led_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                              // led_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [102:0] led_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                       // led_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          led_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                      // id_router_004:sink_ready -> led_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          key_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                // key_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire          key_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                      // key_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire          key_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                              // key_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [102:0] key_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                       // key_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire          key_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                      // id_router_005:sink_ready -> key_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                 // sw_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                       // sw_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                               // sw_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [102:0] sw_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                        // sw_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire          sw_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                       // id_router_006:sink_ready -> sw_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                              // timer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                    // timer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                            // timer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [102:0] timer_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                     // timer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                    // id_router_007:sink_ready -> timer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                           // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [102:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                            // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_008:sink_ready -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire          ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                                  // Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire          ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [102:0] ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                                   // Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire          ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_009:sink_ready -> Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire          ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                                  // Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire          ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire  [102:0] ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                                   // Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire          ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_010:sink_ready -> Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // adc_spi_read_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire          adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                          // adc_spi_read_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire          adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // adc_spi_read_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire  [102:0] adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rp_data;                                           // adc_spi_read_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire          adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_011:sink_ready -> adc_spi_read_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                     // PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire          pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                           // PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire          pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                   // PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire  [102:0] pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data;                                            // PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire          pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                           // id_router_012:sink_ready -> PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                     // PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire          pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                           // PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire          pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                   // PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire  [102:0] pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data;                                            // PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire          pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                           // id_router_013:sink_ready -> PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                       // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	wire  [102:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                                // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                               // id_router_014:sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	wire          encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                                     // encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	wire          encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	wire  [102:0] encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                                      // encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	wire          encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_015:sink_ready -> encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_016:sink_endofpacket
	wire          encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                                     // encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_016:sink_valid
	wire          encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_016:sink_startofpacket
	wire  [102:0] encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                                      // encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_016:sink_data
	wire          encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_016:sink_ready -> encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                              // pio_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_017:sink_endofpacket
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                    // pio_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_017:sink_valid
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                            // pio_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_017:sink_startofpacket
	wire  [102:0] pio_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                     // pio_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_017:sink_data
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                    // id_router_017:sink_ready -> pio_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                             // uart_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_018:sink_endofpacket
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                   // uart_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_018:sink_valid
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                           // uart_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_018:sink_startofpacket
	wire  [102:0] uart_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                    // uart_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_018:sink_data
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                   // id_router_018:sink_ready -> uart_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_019:sink_endofpacket
	wire          ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                                  // Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_019:sink_valid
	wire          ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_019:sink_startofpacket
	wire  [102:0] ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                                   // Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_019:sink_data
	wire          ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_019:sink_ready -> Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_020:sink_endofpacket
	wire          ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                                  // Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_020:sink_valid
	wire          ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_020:sink_startofpacket
	wire  [102:0] ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                                   // Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_020:sink_data
	wire          ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_020:sink_ready -> Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_021:sink_endofpacket
	wire          ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                                  // Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_021:sink_valid
	wire          ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_021:sink_startofpacket
	wire  [102:0] ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                                   // Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_021:sink_data
	wire          ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_021:sink_ready -> Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_022:sink_endofpacket
	wire          ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                                  // Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_022:sink_valid
	wire          ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_022:sink_startofpacket
	wire  [102:0] ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                                   // Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_022:sink_data
	wire          ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_022:sink_ready -> Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                     // PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_023:sink_endofpacket
	wire          pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                           // PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_023:sink_valid
	wire          pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                   // PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_023:sink_startofpacket
	wire  [102:0] pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data;                                            // PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_023:sink_data
	wire          pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                           // id_router_023:sink_ready -> PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                     // PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_024:sink_endofpacket
	wire          pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                           // PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_024:sink_valid
	wire          pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                   // PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_024:sink_startofpacket
	wire  [102:0] pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data;                                            // PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_024:sink_data
	wire          pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                           // id_router_024:sink_ready -> PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                              // pio_1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_025:sink_endofpacket
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                    // pio_1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_025:sink_valid
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                            // pio_1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_025:sink_startofpacket
	wire  [102:0] pio_1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                     // pio_1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_025:sink_data
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                    // id_router_025:sink_ready -> pio_1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          burst_adapter_source0_endofpacket;                                                                              // burst_adapter:source0_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_source0_valid;                                                                                    // burst_adapter:source0_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_source0_startofpacket;                                                                            // burst_adapter:source0_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [84:0] burst_adapter_source0_data;                                                                                     // burst_adapter:source0_data -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_source0_ready;                                                                                    // sdram_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire   [25:0] burst_adapter_source0_channel;                                                                                  // burst_adapter:source0_channel -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rst_controller_reset_out_reset;                                                                                 // rst_controller:reset_out -> [PWM2:csi_I_rst, PWM2_avalon_slave_translator:reset, PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:reset, PWM2_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, PWM3:csi_I_rst, PWM3_avalon_slave_translator:reset, PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:reset, PWM3_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Ultrasound2:reset_n, Ultrasound2_avalon_slave_0_translator:reset, Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Ultrasound3:reset_n, Ultrasound3_avalon_slave_0_translator:reset, Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Ultrasound4:reset_n, Ultrasound4_avalon_slave_0_translator:reset, Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Ultrasound5:reset_n, Ultrasound5_avalon_slave_0_translator:reset, Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, addr_router_001:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_003:reset, crosser:in_reset, crosser_001:out_reset, epcs_flash_controller_0:reset_n, epcs_flash_controller_0_epcs_control_port_translator:reset, epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:reset, epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_003:reset, id_router_018:reset, id_router_019:reset, id_router_020:reset, id_router_021:reset, id_router_022:reset, id_router_023:reset, id_router_024:reset, id_router_025:reset, irq_mapper:reset, nios2_qsys_0:reset_n, nios2_qsys_0_data_master_translator:reset, nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_0_instruction_master_translator:reset, nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_0_jtag_debug_module_translator:reset, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_1:reset_n, pio_1_s1_translator:reset, pio_1_s1_translator_avalon_universal_slave_0_agent:reset, pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_018:reset, rsp_xbar_demux_019:reset, rsp_xbar_demux_020:reset, rsp_xbar_demux_021:reset, rsp_xbar_demux_022:reset, rsp_xbar_demux_023:reset, rsp_xbar_demux_024:reset, rsp_xbar_demux_025:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, uart_0:reset_n, uart_0_s1_translator:reset, uart_0_s1_translator_avalon_universal_slave_0_agent:reset, uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire          rst_controller_001_reset_out_reset;                                                                             // rst_controller_001:reset_out -> [PWM0:csi_I_rst, PWM0_avalon_slave_translator:reset, PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:reset, PWM0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, PWM1:csi_I_rst, PWM1_avalon_slave_translator:reset, PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:reset, PWM1_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Ultrasound0:reset_n, Ultrasound0_avalon_slave_0_translator:reset, Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Ultrasound1:reset_n, Ultrasound1_avalon_slave_0_translator:reset, Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, burst_adapter:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, encoder0:reset_n, encoder0_avalon_slave_0_translator:reset, encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, encoder1:reset_n, encoder1_avalon_slave_0_translator:reset, encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_001:reset, id_router_002:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_012:reset, id_router_013:reset, id_router_014:reset, id_router_015:reset, id_router_016:reset, id_router_017:reset, jtag_uart_0:rst_n, jtag_uart_0_avalon_jtag_slave_translator:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, key:reset_n, key_s1_translator:reset, key_s1_translator_avalon_universal_slave_0_agent:reset, key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, led:reset_n, led_s1_translator:reset, led_s1_translator_avalon_universal_slave_0_agent:reset, led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, onchip_memory2_0:reset, onchip_memory2_0_s1_translator:reset, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:reset, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, performance_counter:reset_n, performance_counter_control_slave_translator:reset, performance_counter_control_slave_translator_avalon_universal_slave_0_agent:reset, performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_0:reset_n, pio_0_s1_translator:reset, pio_0_s1_translator_avalon_universal_slave_0_agent:reset, pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_demux_016:reset, rsp_xbar_demux_017:reset, sdram:reset_n, sdram_s1_translator:reset, sdram_s1_translator_avalon_universal_slave_0_agent:reset, sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sw:reset_n, sw_s1_translator:reset, sw_s1_translator_avalon_universal_slave_0_agent:reset, sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer:reset_n, timer_s1_translator:reset, timer_s1_translator_avalon_universal_slave_0_agent:reset, timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter:reset, width_adapter_001:reset]
	wire          rst_controller_001_reset_out_reset_req;                                                                         // rst_controller_001:reset_req -> onchip_memory2_0:reset_req
	wire          nios2_qsys_0_jtag_debug_module_reset_reset;                                                                     // nios2_qsys_0:jtag_debug_module_resetrequest -> [rst_controller_001:reset_in0, rst_controller_002:reset_in1, rst_controller_003:reset_in1]
	wire          rst_controller_002_reset_out_reset;                                                                             // rst_controller_002:reset_out -> altpll_0:reset
	wire          rst_controller_003_reset_out_reset;                                                                             // rst_controller_003:reset_out -> [adc_spi_read:reset_n, adc_spi_read_slave_translator:reset, adc_spi_read_slave_translator_avalon_universal_slave_0_agent:reset, adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, crosser:out_reset, crosser_001:in_reset, id_router_011:reset, rsp_xbar_demux_011:reset]
	wire          cmd_xbar_demux_src0_endofpacket;                                                                                // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                                      // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                              // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [102:0] cmd_xbar_demux_src0_data;                                                                                       // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [25:0] cmd_xbar_demux_src0_channel;                                                                                    // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire          cmd_xbar_demux_src0_ready;                                                                                      // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire          cmd_xbar_demux_src1_endofpacket;                                                                                // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                                      // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                              // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [102:0] cmd_xbar_demux_src1_data;                                                                                       // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire   [25:0] cmd_xbar_demux_src1_channel;                                                                                    // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire          cmd_xbar_demux_src1_ready;                                                                                      // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire          cmd_xbar_demux_src2_endofpacket;                                                                                // cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire          cmd_xbar_demux_src2_valid;                                                                                      // cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	wire          cmd_xbar_demux_src2_startofpacket;                                                                              // cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [102:0] cmd_xbar_demux_src2_data;                                                                                       // cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	wire   [25:0] cmd_xbar_demux_src2_channel;                                                                                    // cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	wire          cmd_xbar_demux_src2_ready;                                                                                      // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	wire          cmd_xbar_demux_src3_endofpacket;                                                                                // cmd_xbar_demux:src3_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	wire          cmd_xbar_demux_src3_valid;                                                                                      // cmd_xbar_demux:src3_valid -> cmd_xbar_mux_003:sink0_valid
	wire          cmd_xbar_demux_src3_startofpacket;                                                                              // cmd_xbar_demux:src3_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	wire  [102:0] cmd_xbar_demux_src3_data;                                                                                       // cmd_xbar_demux:src3_data -> cmd_xbar_mux_003:sink0_data
	wire   [25:0] cmd_xbar_demux_src3_channel;                                                                                    // cmd_xbar_demux:src3_channel -> cmd_xbar_mux_003:sink0_channel
	wire          cmd_xbar_demux_src3_ready;                                                                                      // cmd_xbar_mux_003:sink0_ready -> cmd_xbar_demux:src3_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                                            // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                                  // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                                          // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src0_data;                                                                                   // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [25:0] cmd_xbar_demux_001_src0_channel;                                                                                // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                                  // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_001_src1_endofpacket;                                                                            // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire          cmd_xbar_demux_001_src1_valid;                                                                                  // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire          cmd_xbar_demux_001_src1_startofpacket;                                                                          // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src1_data;                                                                                   // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire   [25:0] cmd_xbar_demux_001_src1_channel;                                                                                // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire          cmd_xbar_demux_001_src1_ready;                                                                                  // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire          cmd_xbar_demux_001_src2_endofpacket;                                                                            // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire          cmd_xbar_demux_001_src2_valid;                                                                                  // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	wire          cmd_xbar_demux_001_src2_startofpacket;                                                                          // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src2_data;                                                                                   // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	wire   [25:0] cmd_xbar_demux_001_src2_channel;                                                                                // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	wire          cmd_xbar_demux_001_src2_ready;                                                                                  // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	wire          cmd_xbar_demux_001_src3_endofpacket;                                                                            // cmd_xbar_demux_001:src3_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	wire          cmd_xbar_demux_001_src3_valid;                                                                                  // cmd_xbar_demux_001:src3_valid -> cmd_xbar_mux_003:sink1_valid
	wire          cmd_xbar_demux_001_src3_startofpacket;                                                                          // cmd_xbar_demux_001:src3_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src3_data;                                                                                   // cmd_xbar_demux_001:src3_data -> cmd_xbar_mux_003:sink1_data
	wire   [25:0] cmd_xbar_demux_001_src3_channel;                                                                                // cmd_xbar_demux_001:src3_channel -> cmd_xbar_mux_003:sink1_channel
	wire          cmd_xbar_demux_001_src3_ready;                                                                                  // cmd_xbar_mux_003:sink1_ready -> cmd_xbar_demux_001:src3_ready
	wire          cmd_xbar_demux_001_src4_endofpacket;                                                                            // cmd_xbar_demux_001:src4_endofpacket -> led_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src4_valid;                                                                                  // cmd_xbar_demux_001:src4_valid -> led_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src4_startofpacket;                                                                          // cmd_xbar_demux_001:src4_startofpacket -> led_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src4_data;                                                                                   // cmd_xbar_demux_001:src4_data -> led_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [25:0] cmd_xbar_demux_001_src4_channel;                                                                                // cmd_xbar_demux_001:src4_channel -> led_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src5_endofpacket;                                                                            // cmd_xbar_demux_001:src5_endofpacket -> key_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src5_valid;                                                                                  // cmd_xbar_demux_001:src5_valid -> key_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src5_startofpacket;                                                                          // cmd_xbar_demux_001:src5_startofpacket -> key_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src5_data;                                                                                   // cmd_xbar_demux_001:src5_data -> key_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [25:0] cmd_xbar_demux_001_src5_channel;                                                                                // cmd_xbar_demux_001:src5_channel -> key_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src6_endofpacket;                                                                            // cmd_xbar_demux_001:src6_endofpacket -> sw_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src6_valid;                                                                                  // cmd_xbar_demux_001:src6_valid -> sw_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src6_startofpacket;                                                                          // cmd_xbar_demux_001:src6_startofpacket -> sw_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src6_data;                                                                                   // cmd_xbar_demux_001:src6_data -> sw_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [25:0] cmd_xbar_demux_001_src6_channel;                                                                                // cmd_xbar_demux_001:src6_channel -> sw_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src7_endofpacket;                                                                            // cmd_xbar_demux_001:src7_endofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src7_valid;                                                                                  // cmd_xbar_demux_001:src7_valid -> timer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src7_startofpacket;                                                                          // cmd_xbar_demux_001:src7_startofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src7_data;                                                                                   // cmd_xbar_demux_001:src7_data -> timer_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [25:0] cmd_xbar_demux_001_src7_channel;                                                                                // cmd_xbar_demux_001:src7_channel -> timer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src8_endofpacket;                                                                            // cmd_xbar_demux_001:src8_endofpacket -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src8_valid;                                                                                  // cmd_xbar_demux_001:src8_valid -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src8_startofpacket;                                                                          // cmd_xbar_demux_001:src8_startofpacket -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src8_data;                                                                                   // cmd_xbar_demux_001:src8_data -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [25:0] cmd_xbar_demux_001_src8_channel;                                                                                // cmd_xbar_demux_001:src8_channel -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src9_endofpacket;                                                                            // cmd_xbar_demux_001:src9_endofpacket -> Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src9_valid;                                                                                  // cmd_xbar_demux_001:src9_valid -> Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src9_startofpacket;                                                                          // cmd_xbar_demux_001:src9_startofpacket -> Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src9_data;                                                                                   // cmd_xbar_demux_001:src9_data -> Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [25:0] cmd_xbar_demux_001_src9_channel;                                                                                // cmd_xbar_demux_001:src9_channel -> Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src10_endofpacket;                                                                           // cmd_xbar_demux_001:src10_endofpacket -> Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src10_valid;                                                                                 // cmd_xbar_demux_001:src10_valid -> Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src10_startofpacket;                                                                         // cmd_xbar_demux_001:src10_startofpacket -> Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src10_data;                                                                                  // cmd_xbar_demux_001:src10_data -> Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [25:0] cmd_xbar_demux_001_src10_channel;                                                                               // cmd_xbar_demux_001:src10_channel -> Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src12_endofpacket;                                                                           // cmd_xbar_demux_001:src12_endofpacket -> PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src12_valid;                                                                                 // cmd_xbar_demux_001:src12_valid -> PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src12_startofpacket;                                                                         // cmd_xbar_demux_001:src12_startofpacket -> PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src12_data;                                                                                  // cmd_xbar_demux_001:src12_data -> PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [25:0] cmd_xbar_demux_001_src12_channel;                                                                               // cmd_xbar_demux_001:src12_channel -> PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src13_endofpacket;                                                                           // cmd_xbar_demux_001:src13_endofpacket -> PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src13_valid;                                                                                 // cmd_xbar_demux_001:src13_valid -> PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src13_startofpacket;                                                                         // cmd_xbar_demux_001:src13_startofpacket -> PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src13_data;                                                                                  // cmd_xbar_demux_001:src13_data -> PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [25:0] cmd_xbar_demux_001_src13_channel;                                                                               // cmd_xbar_demux_001:src13_channel -> PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src14_endofpacket;                                                                           // cmd_xbar_demux_001:src14_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src14_valid;                                                                                 // cmd_xbar_demux_001:src14_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src14_startofpacket;                                                                         // cmd_xbar_demux_001:src14_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src14_data;                                                                                  // cmd_xbar_demux_001:src14_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [25:0] cmd_xbar_demux_001_src14_channel;                                                                               // cmd_xbar_demux_001:src14_channel -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src15_endofpacket;                                                                           // cmd_xbar_demux_001:src15_endofpacket -> encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src15_valid;                                                                                 // cmd_xbar_demux_001:src15_valid -> encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src15_startofpacket;                                                                         // cmd_xbar_demux_001:src15_startofpacket -> encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src15_data;                                                                                  // cmd_xbar_demux_001:src15_data -> encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [25:0] cmd_xbar_demux_001_src15_channel;                                                                               // cmd_xbar_demux_001:src15_channel -> encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src16_endofpacket;                                                                           // cmd_xbar_demux_001:src16_endofpacket -> encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src16_valid;                                                                                 // cmd_xbar_demux_001:src16_valid -> encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src16_startofpacket;                                                                         // cmd_xbar_demux_001:src16_startofpacket -> encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src16_data;                                                                                  // cmd_xbar_demux_001:src16_data -> encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [25:0] cmd_xbar_demux_001_src16_channel;                                                                               // cmd_xbar_demux_001:src16_channel -> encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src17_endofpacket;                                                                           // cmd_xbar_demux_001:src17_endofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src17_valid;                                                                                 // cmd_xbar_demux_001:src17_valid -> pio_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src17_startofpacket;                                                                         // cmd_xbar_demux_001:src17_startofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src17_data;                                                                                  // cmd_xbar_demux_001:src17_data -> pio_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [25:0] cmd_xbar_demux_001_src17_channel;                                                                               // cmd_xbar_demux_001:src17_channel -> pio_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src18_endofpacket;                                                                           // cmd_xbar_demux_001:src18_endofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src18_valid;                                                                                 // cmd_xbar_demux_001:src18_valid -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src18_startofpacket;                                                                         // cmd_xbar_demux_001:src18_startofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src18_data;                                                                                  // cmd_xbar_demux_001:src18_data -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [25:0] cmd_xbar_demux_001_src18_channel;                                                                               // cmd_xbar_demux_001:src18_channel -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src19_endofpacket;                                                                           // cmd_xbar_demux_001:src19_endofpacket -> Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src19_valid;                                                                                 // cmd_xbar_demux_001:src19_valid -> Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src19_startofpacket;                                                                         // cmd_xbar_demux_001:src19_startofpacket -> Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src19_data;                                                                                  // cmd_xbar_demux_001:src19_data -> Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [25:0] cmd_xbar_demux_001_src19_channel;                                                                               // cmd_xbar_demux_001:src19_channel -> Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src20_endofpacket;                                                                           // cmd_xbar_demux_001:src20_endofpacket -> Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src20_valid;                                                                                 // cmd_xbar_demux_001:src20_valid -> Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src20_startofpacket;                                                                         // cmd_xbar_demux_001:src20_startofpacket -> Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src20_data;                                                                                  // cmd_xbar_demux_001:src20_data -> Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [25:0] cmd_xbar_demux_001_src20_channel;                                                                               // cmd_xbar_demux_001:src20_channel -> Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src21_endofpacket;                                                                           // cmd_xbar_demux_001:src21_endofpacket -> Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src21_valid;                                                                                 // cmd_xbar_demux_001:src21_valid -> Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src21_startofpacket;                                                                         // cmd_xbar_demux_001:src21_startofpacket -> Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src21_data;                                                                                  // cmd_xbar_demux_001:src21_data -> Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [25:0] cmd_xbar_demux_001_src21_channel;                                                                               // cmd_xbar_demux_001:src21_channel -> Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src22_endofpacket;                                                                           // cmd_xbar_demux_001:src22_endofpacket -> Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src22_valid;                                                                                 // cmd_xbar_demux_001:src22_valid -> Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src22_startofpacket;                                                                         // cmd_xbar_demux_001:src22_startofpacket -> Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src22_data;                                                                                  // cmd_xbar_demux_001:src22_data -> Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [25:0] cmd_xbar_demux_001_src22_channel;                                                                               // cmd_xbar_demux_001:src22_channel -> Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src23_endofpacket;                                                                           // cmd_xbar_demux_001:src23_endofpacket -> PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src23_valid;                                                                                 // cmd_xbar_demux_001:src23_valid -> PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src23_startofpacket;                                                                         // cmd_xbar_demux_001:src23_startofpacket -> PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src23_data;                                                                                  // cmd_xbar_demux_001:src23_data -> PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [25:0] cmd_xbar_demux_001_src23_channel;                                                                               // cmd_xbar_demux_001:src23_channel -> PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src24_endofpacket;                                                                           // cmd_xbar_demux_001:src24_endofpacket -> PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src24_valid;                                                                                 // cmd_xbar_demux_001:src24_valid -> PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src24_startofpacket;                                                                         // cmd_xbar_demux_001:src24_startofpacket -> PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src24_data;                                                                                  // cmd_xbar_demux_001:src24_data -> PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [25:0] cmd_xbar_demux_001_src24_channel;                                                                               // cmd_xbar_demux_001:src24_channel -> PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src25_endofpacket;                                                                           // cmd_xbar_demux_001:src25_endofpacket -> pio_1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src25_valid;                                                                                 // cmd_xbar_demux_001:src25_valid -> pio_1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src25_startofpacket;                                                                         // cmd_xbar_demux_001:src25_startofpacket -> pio_1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src25_data;                                                                                  // cmd_xbar_demux_001:src25_data -> pio_1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [25:0] cmd_xbar_demux_001_src25_channel;                                                                               // cmd_xbar_demux_001:src25_channel -> pio_1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rsp_xbar_demux_src0_endofpacket;                                                                                // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                                      // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                              // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [102:0] rsp_xbar_demux_src0_data;                                                                                       // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [25:0] rsp_xbar_demux_src0_channel;                                                                                    // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                                      // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_src1_endofpacket;                                                                                // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                                                      // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                                                              // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [102:0] rsp_xbar_demux_src1_data;                                                                                       // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire   [25:0] rsp_xbar_demux_src1_channel;                                                                                    // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire          rsp_xbar_demux_src1_ready;                                                                                      // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                                            // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                                  // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                                          // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [102:0] rsp_xbar_demux_001_src0_data;                                                                                   // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [25:0] rsp_xbar_demux_001_src0_channel;                                                                                // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                                  // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_001_src1_endofpacket;                                                                            // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire          rsp_xbar_demux_001_src1_valid;                                                                                  // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire          rsp_xbar_demux_001_src1_startofpacket;                                                                          // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [102:0] rsp_xbar_demux_001_src1_data;                                                                                   // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire   [25:0] rsp_xbar_demux_001_src1_channel;                                                                                // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire          rsp_xbar_demux_001_src1_ready;                                                                                  // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                                            // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                                  // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                                          // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [102:0] rsp_xbar_demux_002_src0_data;                                                                                   // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire   [25:0] rsp_xbar_demux_002_src0_channel;                                                                                // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                                  // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_002_src1_endofpacket;                                                                            // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire          rsp_xbar_demux_002_src1_valid;                                                                                  // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	wire          rsp_xbar_demux_002_src1_startofpacket;                                                                          // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [102:0] rsp_xbar_demux_002_src1_data;                                                                                   // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	wire   [25:0] rsp_xbar_demux_002_src1_channel;                                                                                // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	wire          rsp_xbar_demux_002_src1_ready;                                                                                  // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                                            // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                                  // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                                          // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire  [102:0] rsp_xbar_demux_003_src0_data;                                                                                   // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	wire   [25:0] rsp_xbar_demux_003_src0_channel;                                                                                // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                                  // rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_003_src1_endofpacket;                                                                            // rsp_xbar_demux_003:src1_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire          rsp_xbar_demux_003_src1_valid;                                                                                  // rsp_xbar_demux_003:src1_valid -> rsp_xbar_mux_001:sink3_valid
	wire          rsp_xbar_demux_003_src1_startofpacket;                                                                          // rsp_xbar_demux_003:src1_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [102:0] rsp_xbar_demux_003_src1_data;                                                                                   // rsp_xbar_demux_003:src1_data -> rsp_xbar_mux_001:sink3_data
	wire   [25:0] rsp_xbar_demux_003_src1_channel;                                                                                // rsp_xbar_demux_003:src1_channel -> rsp_xbar_mux_001:sink3_channel
	wire          rsp_xbar_demux_003_src1_ready;                                                                                  // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src1_ready
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                                            // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                                  // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink4_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                                          // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [102:0] rsp_xbar_demux_004_src0_data;                                                                                   // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink4_data
	wire   [25:0] rsp_xbar_demux_004_src0_channel;                                                                                // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink4_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                                  // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                                            // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                                  // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                                          // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [102:0] rsp_xbar_demux_005_src0_data;                                                                                   // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	wire   [25:0] rsp_xbar_demux_005_src0_channel;                                                                                // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	wire          rsp_xbar_demux_005_src0_ready;                                                                                  // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire          rsp_xbar_demux_006_src0_endofpacket;                                                                            // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire          rsp_xbar_demux_006_src0_valid;                                                                                  // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	wire          rsp_xbar_demux_006_src0_startofpacket;                                                                          // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [102:0] rsp_xbar_demux_006_src0_data;                                                                                   // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	wire   [25:0] rsp_xbar_demux_006_src0_channel;                                                                                // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	wire          rsp_xbar_demux_006_src0_ready;                                                                                  // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire          rsp_xbar_demux_007_src0_endofpacket;                                                                            // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire          rsp_xbar_demux_007_src0_valid;                                                                                  // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	wire          rsp_xbar_demux_007_src0_startofpacket;                                                                          // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [102:0] rsp_xbar_demux_007_src0_data;                                                                                   // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	wire   [25:0] rsp_xbar_demux_007_src0_channel;                                                                                // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	wire          rsp_xbar_demux_007_src0_ready;                                                                                  // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire          rsp_xbar_demux_008_src0_endofpacket;                                                                            // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire          rsp_xbar_demux_008_src0_valid;                                                                                  // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	wire          rsp_xbar_demux_008_src0_startofpacket;                                                                          // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [102:0] rsp_xbar_demux_008_src0_data;                                                                                   // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	wire   [25:0] rsp_xbar_demux_008_src0_channel;                                                                                // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	wire          rsp_xbar_demux_008_src0_ready;                                                                                  // rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire          rsp_xbar_demux_009_src0_endofpacket;                                                                            // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	wire          rsp_xbar_demux_009_src0_valid;                                                                                  // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_001:sink9_valid
	wire          rsp_xbar_demux_009_src0_startofpacket;                                                                          // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	wire  [102:0] rsp_xbar_demux_009_src0_data;                                                                                   // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_001:sink9_data
	wire   [25:0] rsp_xbar_demux_009_src0_channel;                                                                                // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_001:sink9_channel
	wire          rsp_xbar_demux_009_src0_ready;                                                                                  // rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src0_ready
	wire          rsp_xbar_demux_010_src0_endofpacket;                                                                            // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	wire          rsp_xbar_demux_010_src0_valid;                                                                                  // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_001:sink10_valid
	wire          rsp_xbar_demux_010_src0_startofpacket;                                                                          // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	wire  [102:0] rsp_xbar_demux_010_src0_data;                                                                                   // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_001:sink10_data
	wire   [25:0] rsp_xbar_demux_010_src0_channel;                                                                                // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_001:sink10_channel
	wire          rsp_xbar_demux_010_src0_ready;                                                                                  // rsp_xbar_mux_001:sink10_ready -> rsp_xbar_demux_010:src0_ready
	wire          rsp_xbar_demux_012_src0_endofpacket;                                                                            // rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux_001:sink12_endofpacket
	wire          rsp_xbar_demux_012_src0_valid;                                                                                  // rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux_001:sink12_valid
	wire          rsp_xbar_demux_012_src0_startofpacket;                                                                          // rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux_001:sink12_startofpacket
	wire  [102:0] rsp_xbar_demux_012_src0_data;                                                                                   // rsp_xbar_demux_012:src0_data -> rsp_xbar_mux_001:sink12_data
	wire   [25:0] rsp_xbar_demux_012_src0_channel;                                                                                // rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux_001:sink12_channel
	wire          rsp_xbar_demux_012_src0_ready;                                                                                  // rsp_xbar_mux_001:sink12_ready -> rsp_xbar_demux_012:src0_ready
	wire          rsp_xbar_demux_013_src0_endofpacket;                                                                            // rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux_001:sink13_endofpacket
	wire          rsp_xbar_demux_013_src0_valid;                                                                                  // rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux_001:sink13_valid
	wire          rsp_xbar_demux_013_src0_startofpacket;                                                                          // rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux_001:sink13_startofpacket
	wire  [102:0] rsp_xbar_demux_013_src0_data;                                                                                   // rsp_xbar_demux_013:src0_data -> rsp_xbar_mux_001:sink13_data
	wire   [25:0] rsp_xbar_demux_013_src0_channel;                                                                                // rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux_001:sink13_channel
	wire          rsp_xbar_demux_013_src0_ready;                                                                                  // rsp_xbar_mux_001:sink13_ready -> rsp_xbar_demux_013:src0_ready
	wire          rsp_xbar_demux_014_src0_endofpacket;                                                                            // rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux_001:sink14_endofpacket
	wire          rsp_xbar_demux_014_src0_valid;                                                                                  // rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux_001:sink14_valid
	wire          rsp_xbar_demux_014_src0_startofpacket;                                                                          // rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux_001:sink14_startofpacket
	wire  [102:0] rsp_xbar_demux_014_src0_data;                                                                                   // rsp_xbar_demux_014:src0_data -> rsp_xbar_mux_001:sink14_data
	wire   [25:0] rsp_xbar_demux_014_src0_channel;                                                                                // rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux_001:sink14_channel
	wire          rsp_xbar_demux_014_src0_ready;                                                                                  // rsp_xbar_mux_001:sink14_ready -> rsp_xbar_demux_014:src0_ready
	wire          rsp_xbar_demux_015_src0_endofpacket;                                                                            // rsp_xbar_demux_015:src0_endofpacket -> rsp_xbar_mux_001:sink15_endofpacket
	wire          rsp_xbar_demux_015_src0_valid;                                                                                  // rsp_xbar_demux_015:src0_valid -> rsp_xbar_mux_001:sink15_valid
	wire          rsp_xbar_demux_015_src0_startofpacket;                                                                          // rsp_xbar_demux_015:src0_startofpacket -> rsp_xbar_mux_001:sink15_startofpacket
	wire  [102:0] rsp_xbar_demux_015_src0_data;                                                                                   // rsp_xbar_demux_015:src0_data -> rsp_xbar_mux_001:sink15_data
	wire   [25:0] rsp_xbar_demux_015_src0_channel;                                                                                // rsp_xbar_demux_015:src0_channel -> rsp_xbar_mux_001:sink15_channel
	wire          rsp_xbar_demux_015_src0_ready;                                                                                  // rsp_xbar_mux_001:sink15_ready -> rsp_xbar_demux_015:src0_ready
	wire          rsp_xbar_demux_016_src0_endofpacket;                                                                            // rsp_xbar_demux_016:src0_endofpacket -> rsp_xbar_mux_001:sink16_endofpacket
	wire          rsp_xbar_demux_016_src0_valid;                                                                                  // rsp_xbar_demux_016:src0_valid -> rsp_xbar_mux_001:sink16_valid
	wire          rsp_xbar_demux_016_src0_startofpacket;                                                                          // rsp_xbar_demux_016:src0_startofpacket -> rsp_xbar_mux_001:sink16_startofpacket
	wire  [102:0] rsp_xbar_demux_016_src0_data;                                                                                   // rsp_xbar_demux_016:src0_data -> rsp_xbar_mux_001:sink16_data
	wire   [25:0] rsp_xbar_demux_016_src0_channel;                                                                                // rsp_xbar_demux_016:src0_channel -> rsp_xbar_mux_001:sink16_channel
	wire          rsp_xbar_demux_016_src0_ready;                                                                                  // rsp_xbar_mux_001:sink16_ready -> rsp_xbar_demux_016:src0_ready
	wire          rsp_xbar_demux_017_src0_endofpacket;                                                                            // rsp_xbar_demux_017:src0_endofpacket -> rsp_xbar_mux_001:sink17_endofpacket
	wire          rsp_xbar_demux_017_src0_valid;                                                                                  // rsp_xbar_demux_017:src0_valid -> rsp_xbar_mux_001:sink17_valid
	wire          rsp_xbar_demux_017_src0_startofpacket;                                                                          // rsp_xbar_demux_017:src0_startofpacket -> rsp_xbar_mux_001:sink17_startofpacket
	wire  [102:0] rsp_xbar_demux_017_src0_data;                                                                                   // rsp_xbar_demux_017:src0_data -> rsp_xbar_mux_001:sink17_data
	wire   [25:0] rsp_xbar_demux_017_src0_channel;                                                                                // rsp_xbar_demux_017:src0_channel -> rsp_xbar_mux_001:sink17_channel
	wire          rsp_xbar_demux_017_src0_ready;                                                                                  // rsp_xbar_mux_001:sink17_ready -> rsp_xbar_demux_017:src0_ready
	wire          rsp_xbar_demux_018_src0_endofpacket;                                                                            // rsp_xbar_demux_018:src0_endofpacket -> rsp_xbar_mux_001:sink18_endofpacket
	wire          rsp_xbar_demux_018_src0_valid;                                                                                  // rsp_xbar_demux_018:src0_valid -> rsp_xbar_mux_001:sink18_valid
	wire          rsp_xbar_demux_018_src0_startofpacket;                                                                          // rsp_xbar_demux_018:src0_startofpacket -> rsp_xbar_mux_001:sink18_startofpacket
	wire  [102:0] rsp_xbar_demux_018_src0_data;                                                                                   // rsp_xbar_demux_018:src0_data -> rsp_xbar_mux_001:sink18_data
	wire   [25:0] rsp_xbar_demux_018_src0_channel;                                                                                // rsp_xbar_demux_018:src0_channel -> rsp_xbar_mux_001:sink18_channel
	wire          rsp_xbar_demux_018_src0_ready;                                                                                  // rsp_xbar_mux_001:sink18_ready -> rsp_xbar_demux_018:src0_ready
	wire          rsp_xbar_demux_019_src0_endofpacket;                                                                            // rsp_xbar_demux_019:src0_endofpacket -> rsp_xbar_mux_001:sink19_endofpacket
	wire          rsp_xbar_demux_019_src0_valid;                                                                                  // rsp_xbar_demux_019:src0_valid -> rsp_xbar_mux_001:sink19_valid
	wire          rsp_xbar_demux_019_src0_startofpacket;                                                                          // rsp_xbar_demux_019:src0_startofpacket -> rsp_xbar_mux_001:sink19_startofpacket
	wire  [102:0] rsp_xbar_demux_019_src0_data;                                                                                   // rsp_xbar_demux_019:src0_data -> rsp_xbar_mux_001:sink19_data
	wire   [25:0] rsp_xbar_demux_019_src0_channel;                                                                                // rsp_xbar_demux_019:src0_channel -> rsp_xbar_mux_001:sink19_channel
	wire          rsp_xbar_demux_019_src0_ready;                                                                                  // rsp_xbar_mux_001:sink19_ready -> rsp_xbar_demux_019:src0_ready
	wire          rsp_xbar_demux_020_src0_endofpacket;                                                                            // rsp_xbar_demux_020:src0_endofpacket -> rsp_xbar_mux_001:sink20_endofpacket
	wire          rsp_xbar_demux_020_src0_valid;                                                                                  // rsp_xbar_demux_020:src0_valid -> rsp_xbar_mux_001:sink20_valid
	wire          rsp_xbar_demux_020_src0_startofpacket;                                                                          // rsp_xbar_demux_020:src0_startofpacket -> rsp_xbar_mux_001:sink20_startofpacket
	wire  [102:0] rsp_xbar_demux_020_src0_data;                                                                                   // rsp_xbar_demux_020:src0_data -> rsp_xbar_mux_001:sink20_data
	wire   [25:0] rsp_xbar_demux_020_src0_channel;                                                                                // rsp_xbar_demux_020:src0_channel -> rsp_xbar_mux_001:sink20_channel
	wire          rsp_xbar_demux_020_src0_ready;                                                                                  // rsp_xbar_mux_001:sink20_ready -> rsp_xbar_demux_020:src0_ready
	wire          rsp_xbar_demux_021_src0_endofpacket;                                                                            // rsp_xbar_demux_021:src0_endofpacket -> rsp_xbar_mux_001:sink21_endofpacket
	wire          rsp_xbar_demux_021_src0_valid;                                                                                  // rsp_xbar_demux_021:src0_valid -> rsp_xbar_mux_001:sink21_valid
	wire          rsp_xbar_demux_021_src0_startofpacket;                                                                          // rsp_xbar_demux_021:src0_startofpacket -> rsp_xbar_mux_001:sink21_startofpacket
	wire  [102:0] rsp_xbar_demux_021_src0_data;                                                                                   // rsp_xbar_demux_021:src0_data -> rsp_xbar_mux_001:sink21_data
	wire   [25:0] rsp_xbar_demux_021_src0_channel;                                                                                // rsp_xbar_demux_021:src0_channel -> rsp_xbar_mux_001:sink21_channel
	wire          rsp_xbar_demux_021_src0_ready;                                                                                  // rsp_xbar_mux_001:sink21_ready -> rsp_xbar_demux_021:src0_ready
	wire          rsp_xbar_demux_022_src0_endofpacket;                                                                            // rsp_xbar_demux_022:src0_endofpacket -> rsp_xbar_mux_001:sink22_endofpacket
	wire          rsp_xbar_demux_022_src0_valid;                                                                                  // rsp_xbar_demux_022:src0_valid -> rsp_xbar_mux_001:sink22_valid
	wire          rsp_xbar_demux_022_src0_startofpacket;                                                                          // rsp_xbar_demux_022:src0_startofpacket -> rsp_xbar_mux_001:sink22_startofpacket
	wire  [102:0] rsp_xbar_demux_022_src0_data;                                                                                   // rsp_xbar_demux_022:src0_data -> rsp_xbar_mux_001:sink22_data
	wire   [25:0] rsp_xbar_demux_022_src0_channel;                                                                                // rsp_xbar_demux_022:src0_channel -> rsp_xbar_mux_001:sink22_channel
	wire          rsp_xbar_demux_022_src0_ready;                                                                                  // rsp_xbar_mux_001:sink22_ready -> rsp_xbar_demux_022:src0_ready
	wire          rsp_xbar_demux_023_src0_endofpacket;                                                                            // rsp_xbar_demux_023:src0_endofpacket -> rsp_xbar_mux_001:sink23_endofpacket
	wire          rsp_xbar_demux_023_src0_valid;                                                                                  // rsp_xbar_demux_023:src0_valid -> rsp_xbar_mux_001:sink23_valid
	wire          rsp_xbar_demux_023_src0_startofpacket;                                                                          // rsp_xbar_demux_023:src0_startofpacket -> rsp_xbar_mux_001:sink23_startofpacket
	wire  [102:0] rsp_xbar_demux_023_src0_data;                                                                                   // rsp_xbar_demux_023:src0_data -> rsp_xbar_mux_001:sink23_data
	wire   [25:0] rsp_xbar_demux_023_src0_channel;                                                                                // rsp_xbar_demux_023:src0_channel -> rsp_xbar_mux_001:sink23_channel
	wire          rsp_xbar_demux_023_src0_ready;                                                                                  // rsp_xbar_mux_001:sink23_ready -> rsp_xbar_demux_023:src0_ready
	wire          rsp_xbar_demux_024_src0_endofpacket;                                                                            // rsp_xbar_demux_024:src0_endofpacket -> rsp_xbar_mux_001:sink24_endofpacket
	wire          rsp_xbar_demux_024_src0_valid;                                                                                  // rsp_xbar_demux_024:src0_valid -> rsp_xbar_mux_001:sink24_valid
	wire          rsp_xbar_demux_024_src0_startofpacket;                                                                          // rsp_xbar_demux_024:src0_startofpacket -> rsp_xbar_mux_001:sink24_startofpacket
	wire  [102:0] rsp_xbar_demux_024_src0_data;                                                                                   // rsp_xbar_demux_024:src0_data -> rsp_xbar_mux_001:sink24_data
	wire   [25:0] rsp_xbar_demux_024_src0_channel;                                                                                // rsp_xbar_demux_024:src0_channel -> rsp_xbar_mux_001:sink24_channel
	wire          rsp_xbar_demux_024_src0_ready;                                                                                  // rsp_xbar_mux_001:sink24_ready -> rsp_xbar_demux_024:src0_ready
	wire          rsp_xbar_demux_025_src0_endofpacket;                                                                            // rsp_xbar_demux_025:src0_endofpacket -> rsp_xbar_mux_001:sink25_endofpacket
	wire          rsp_xbar_demux_025_src0_valid;                                                                                  // rsp_xbar_demux_025:src0_valid -> rsp_xbar_mux_001:sink25_valid
	wire          rsp_xbar_demux_025_src0_startofpacket;                                                                          // rsp_xbar_demux_025:src0_startofpacket -> rsp_xbar_mux_001:sink25_startofpacket
	wire  [102:0] rsp_xbar_demux_025_src0_data;                                                                                   // rsp_xbar_demux_025:src0_data -> rsp_xbar_mux_001:sink25_data
	wire   [25:0] rsp_xbar_demux_025_src0_channel;                                                                                // rsp_xbar_demux_025:src0_channel -> rsp_xbar_mux_001:sink25_channel
	wire          rsp_xbar_demux_025_src0_ready;                                                                                  // rsp_xbar_mux_001:sink25_ready -> rsp_xbar_demux_025:src0_ready
	wire          addr_router_src_endofpacket;                                                                                    // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          addr_router_src_valid;                                                                                          // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire          addr_router_src_startofpacket;                                                                                  // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [102:0] addr_router_src_data;                                                                                           // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire   [25:0] addr_router_src_channel;                                                                                        // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire          addr_router_src_ready;                                                                                          // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                                   // rsp_xbar_mux:src_endofpacket -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                                         // rsp_xbar_mux:src_valid -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                                 // rsp_xbar_mux:src_startofpacket -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [102:0] rsp_xbar_mux_src_data;                                                                                          // rsp_xbar_mux:src_data -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [25:0] rsp_xbar_mux_src_channel;                                                                                       // rsp_xbar_mux:src_channel -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_src_ready;                                                                                         // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	wire          addr_router_001_src_endofpacket;                                                                                // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          addr_router_001_src_valid;                                                                                      // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire          addr_router_001_src_startofpacket;                                                                              // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [102:0] addr_router_001_src_data;                                                                                       // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire   [25:0] addr_router_001_src_channel;                                                                                    // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire          addr_router_001_src_ready;                                                                                      // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire          rsp_xbar_mux_001_src_endofpacket;                                                                               // rsp_xbar_mux_001:src_endofpacket -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_001_src_valid;                                                                                     // rsp_xbar_mux_001:src_valid -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_001_src_startofpacket;                                                                             // rsp_xbar_mux_001:src_startofpacket -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [102:0] rsp_xbar_mux_001_src_data;                                                                                      // rsp_xbar_mux_001:src_data -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [25:0] rsp_xbar_mux_001_src_channel;                                                                                   // rsp_xbar_mux_001:src_channel -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_001_src_ready;                                                                                     // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	wire          cmd_xbar_mux_src_endofpacket;                                                                                   // cmd_xbar_mux:src_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                                                         // cmd_xbar_mux:src_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                                                 // cmd_xbar_mux:src_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_mux_src_data;                                                                                          // cmd_xbar_mux:src_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [25:0] cmd_xbar_mux_src_channel;                                                                                       // cmd_xbar_mux:src_channel -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_src_ready;                                                                                         // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire          id_router_src_endofpacket;                                                                                      // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                                            // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                                    // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [102:0] id_router_src_data;                                                                                             // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [25:0] id_router_src_channel;                                                                                          // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                                            // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_mux_002_src_endofpacket;                                                                               // cmd_xbar_mux_002:src_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_002_src_valid;                                                                                     // cmd_xbar_mux_002:src_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_002_src_startofpacket;                                                                             // cmd_xbar_mux_002:src_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_mux_002_src_data;                                                                                      // cmd_xbar_mux_002:src_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [25:0] cmd_xbar_mux_002_src_channel;                                                                                   // cmd_xbar_mux_002:src_channel -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_002_src_ready;                                                                                     // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_002:src_ready
	wire          id_router_002_src_endofpacket;                                                                                  // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                                        // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                                                // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [102:0] id_router_002_src_data;                                                                                         // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire   [25:0] id_router_002_src_channel;                                                                                      // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                                        // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire          cmd_xbar_mux_003_src_endofpacket;                                                                               // cmd_xbar_mux_003:src_endofpacket -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_003_src_valid;                                                                                     // cmd_xbar_mux_003:src_valid -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_003_src_startofpacket;                                                                             // cmd_xbar_mux_003:src_startofpacket -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_mux_003_src_data;                                                                                      // cmd_xbar_mux_003:src_data -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_data
	wire   [25:0] cmd_xbar_mux_003_src_channel;                                                                                   // cmd_xbar_mux_003:src_channel -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_003_src_ready;                                                                                     // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_003:src_ready
	wire          id_router_003_src_endofpacket;                                                                                  // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                                        // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                                                // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [102:0] id_router_003_src_data;                                                                                         // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [25:0] id_router_003_src_channel;                                                                                      // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                                        // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          cmd_xbar_demux_001_src4_ready;                                                                                  // led_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	wire          id_router_004_src_endofpacket;                                                                                  // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          id_router_004_src_valid;                                                                                        // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire          id_router_004_src_startofpacket;                                                                                // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [102:0] id_router_004_src_data;                                                                                         // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire   [25:0] id_router_004_src_channel;                                                                                      // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire          id_router_004_src_ready;                                                                                        // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire          cmd_xbar_demux_001_src5_ready;                                                                                  // key_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	wire          id_router_005_src_endofpacket;                                                                                  // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          id_router_005_src_valid;                                                                                        // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire          id_router_005_src_startofpacket;                                                                                // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [102:0] id_router_005_src_data;                                                                                         // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [25:0] id_router_005_src_channel;                                                                                      // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire          id_router_005_src_ready;                                                                                        // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire          cmd_xbar_demux_001_src6_ready;                                                                                  // sw_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	wire          id_router_006_src_endofpacket;                                                                                  // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire          id_router_006_src_valid;                                                                                        // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire          id_router_006_src_startofpacket;                                                                                // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [102:0] id_router_006_src_data;                                                                                         // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire   [25:0] id_router_006_src_channel;                                                                                      // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire          id_router_006_src_ready;                                                                                        // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire          cmd_xbar_demux_001_src7_ready;                                                                                  // timer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	wire          id_router_007_src_endofpacket;                                                                                  // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire          id_router_007_src_valid;                                                                                        // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire          id_router_007_src_startofpacket;                                                                                // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [102:0] id_router_007_src_data;                                                                                         // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire   [25:0] id_router_007_src_channel;                                                                                      // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire          id_router_007_src_ready;                                                                                        // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire          cmd_xbar_demux_001_src8_ready;                                                                                  // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src8_ready
	wire          id_router_008_src_endofpacket;                                                                                  // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire          id_router_008_src_valid;                                                                                        // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire          id_router_008_src_startofpacket;                                                                                // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [102:0] id_router_008_src_data;                                                                                         // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire   [25:0] id_router_008_src_channel;                                                                                      // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire          id_router_008_src_ready;                                                                                        // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire          cmd_xbar_demux_001_src9_ready;                                                                                  // Ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src9_ready
	wire          id_router_009_src_endofpacket;                                                                                  // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire          id_router_009_src_valid;                                                                                        // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire          id_router_009_src_startofpacket;                                                                                // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [102:0] id_router_009_src_data;                                                                                         // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire   [25:0] id_router_009_src_channel;                                                                                      // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire          id_router_009_src_ready;                                                                                        // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire          cmd_xbar_demux_001_src10_ready;                                                                                 // Ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src10_ready
	wire          id_router_010_src_endofpacket;                                                                                  // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire          id_router_010_src_valid;                                                                                        // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire          id_router_010_src_startofpacket;                                                                                // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [102:0] id_router_010_src_data;                                                                                         // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire   [25:0] id_router_010_src_channel;                                                                                      // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire          id_router_010_src_ready;                                                                                        // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire          crosser_out_ready;                                                                                              // adc_spi_read_slave_translator_avalon_universal_slave_0_agent:cp_ready -> crosser:out_ready
	wire          id_router_011_src_endofpacket;                                                                                  // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire          id_router_011_src_valid;                                                                                        // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire          id_router_011_src_startofpacket;                                                                                // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire  [102:0] id_router_011_src_data;                                                                                         // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire   [25:0] id_router_011_src_channel;                                                                                      // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire          id_router_011_src_ready;                                                                                        // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire          cmd_xbar_demux_001_src12_ready;                                                                                 // PWM0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src12_ready
	wire          id_router_012_src_endofpacket;                                                                                  // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire          id_router_012_src_valid;                                                                                        // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire          id_router_012_src_startofpacket;                                                                                // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire  [102:0] id_router_012_src_data;                                                                                         // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire   [25:0] id_router_012_src_channel;                                                                                      // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire          id_router_012_src_ready;                                                                                        // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire          cmd_xbar_demux_001_src13_ready;                                                                                 // PWM1_avalon_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src13_ready
	wire          id_router_013_src_endofpacket;                                                                                  // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire          id_router_013_src_valid;                                                                                        // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire          id_router_013_src_startofpacket;                                                                                // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire  [102:0] id_router_013_src_data;                                                                                         // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire   [25:0] id_router_013_src_channel;                                                                                      // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire          id_router_013_src_ready;                                                                                        // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire          cmd_xbar_demux_001_src14_ready;                                                                                 // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src14_ready
	wire          id_router_014_src_endofpacket;                                                                                  // id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	wire          id_router_014_src_valid;                                                                                        // id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	wire          id_router_014_src_startofpacket;                                                                                // id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	wire  [102:0] id_router_014_src_data;                                                                                         // id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	wire   [25:0] id_router_014_src_channel;                                                                                      // id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	wire          id_router_014_src_ready;                                                                                        // rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	wire          cmd_xbar_demux_001_src15_ready;                                                                                 // encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src15_ready
	wire          id_router_015_src_endofpacket;                                                                                  // id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	wire          id_router_015_src_valid;                                                                                        // id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	wire          id_router_015_src_startofpacket;                                                                                // id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	wire  [102:0] id_router_015_src_data;                                                                                         // id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	wire   [25:0] id_router_015_src_channel;                                                                                      // id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	wire          id_router_015_src_ready;                                                                                        // rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	wire          cmd_xbar_demux_001_src16_ready;                                                                                 // encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src16_ready
	wire          id_router_016_src_endofpacket;                                                                                  // id_router_016:src_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	wire          id_router_016_src_valid;                                                                                        // id_router_016:src_valid -> rsp_xbar_demux_016:sink_valid
	wire          id_router_016_src_startofpacket;                                                                                // id_router_016:src_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	wire  [102:0] id_router_016_src_data;                                                                                         // id_router_016:src_data -> rsp_xbar_demux_016:sink_data
	wire   [25:0] id_router_016_src_channel;                                                                                      // id_router_016:src_channel -> rsp_xbar_demux_016:sink_channel
	wire          id_router_016_src_ready;                                                                                        // rsp_xbar_demux_016:sink_ready -> id_router_016:src_ready
	wire          cmd_xbar_demux_001_src17_ready;                                                                                 // pio_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src17_ready
	wire          id_router_017_src_endofpacket;                                                                                  // id_router_017:src_endofpacket -> rsp_xbar_demux_017:sink_endofpacket
	wire          id_router_017_src_valid;                                                                                        // id_router_017:src_valid -> rsp_xbar_demux_017:sink_valid
	wire          id_router_017_src_startofpacket;                                                                                // id_router_017:src_startofpacket -> rsp_xbar_demux_017:sink_startofpacket
	wire  [102:0] id_router_017_src_data;                                                                                         // id_router_017:src_data -> rsp_xbar_demux_017:sink_data
	wire   [25:0] id_router_017_src_channel;                                                                                      // id_router_017:src_channel -> rsp_xbar_demux_017:sink_channel
	wire          id_router_017_src_ready;                                                                                        // rsp_xbar_demux_017:sink_ready -> id_router_017:src_ready
	wire          cmd_xbar_demux_001_src18_ready;                                                                                 // uart_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src18_ready
	wire          id_router_018_src_endofpacket;                                                                                  // id_router_018:src_endofpacket -> rsp_xbar_demux_018:sink_endofpacket
	wire          id_router_018_src_valid;                                                                                        // id_router_018:src_valid -> rsp_xbar_demux_018:sink_valid
	wire          id_router_018_src_startofpacket;                                                                                // id_router_018:src_startofpacket -> rsp_xbar_demux_018:sink_startofpacket
	wire  [102:0] id_router_018_src_data;                                                                                         // id_router_018:src_data -> rsp_xbar_demux_018:sink_data
	wire   [25:0] id_router_018_src_channel;                                                                                      // id_router_018:src_channel -> rsp_xbar_demux_018:sink_channel
	wire          id_router_018_src_ready;                                                                                        // rsp_xbar_demux_018:sink_ready -> id_router_018:src_ready
	wire          cmd_xbar_demux_001_src19_ready;                                                                                 // Ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src19_ready
	wire          id_router_019_src_endofpacket;                                                                                  // id_router_019:src_endofpacket -> rsp_xbar_demux_019:sink_endofpacket
	wire          id_router_019_src_valid;                                                                                        // id_router_019:src_valid -> rsp_xbar_demux_019:sink_valid
	wire          id_router_019_src_startofpacket;                                                                                // id_router_019:src_startofpacket -> rsp_xbar_demux_019:sink_startofpacket
	wire  [102:0] id_router_019_src_data;                                                                                         // id_router_019:src_data -> rsp_xbar_demux_019:sink_data
	wire   [25:0] id_router_019_src_channel;                                                                                      // id_router_019:src_channel -> rsp_xbar_demux_019:sink_channel
	wire          id_router_019_src_ready;                                                                                        // rsp_xbar_demux_019:sink_ready -> id_router_019:src_ready
	wire          cmd_xbar_demux_001_src20_ready;                                                                                 // Ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src20_ready
	wire          id_router_020_src_endofpacket;                                                                                  // id_router_020:src_endofpacket -> rsp_xbar_demux_020:sink_endofpacket
	wire          id_router_020_src_valid;                                                                                        // id_router_020:src_valid -> rsp_xbar_demux_020:sink_valid
	wire          id_router_020_src_startofpacket;                                                                                // id_router_020:src_startofpacket -> rsp_xbar_demux_020:sink_startofpacket
	wire  [102:0] id_router_020_src_data;                                                                                         // id_router_020:src_data -> rsp_xbar_demux_020:sink_data
	wire   [25:0] id_router_020_src_channel;                                                                                      // id_router_020:src_channel -> rsp_xbar_demux_020:sink_channel
	wire          id_router_020_src_ready;                                                                                        // rsp_xbar_demux_020:sink_ready -> id_router_020:src_ready
	wire          cmd_xbar_demux_001_src21_ready;                                                                                 // Ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src21_ready
	wire          id_router_021_src_endofpacket;                                                                                  // id_router_021:src_endofpacket -> rsp_xbar_demux_021:sink_endofpacket
	wire          id_router_021_src_valid;                                                                                        // id_router_021:src_valid -> rsp_xbar_demux_021:sink_valid
	wire          id_router_021_src_startofpacket;                                                                                // id_router_021:src_startofpacket -> rsp_xbar_demux_021:sink_startofpacket
	wire  [102:0] id_router_021_src_data;                                                                                         // id_router_021:src_data -> rsp_xbar_demux_021:sink_data
	wire   [25:0] id_router_021_src_channel;                                                                                      // id_router_021:src_channel -> rsp_xbar_demux_021:sink_channel
	wire          id_router_021_src_ready;                                                                                        // rsp_xbar_demux_021:sink_ready -> id_router_021:src_ready
	wire          cmd_xbar_demux_001_src22_ready;                                                                                 // Ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src22_ready
	wire          id_router_022_src_endofpacket;                                                                                  // id_router_022:src_endofpacket -> rsp_xbar_demux_022:sink_endofpacket
	wire          id_router_022_src_valid;                                                                                        // id_router_022:src_valid -> rsp_xbar_demux_022:sink_valid
	wire          id_router_022_src_startofpacket;                                                                                // id_router_022:src_startofpacket -> rsp_xbar_demux_022:sink_startofpacket
	wire  [102:0] id_router_022_src_data;                                                                                         // id_router_022:src_data -> rsp_xbar_demux_022:sink_data
	wire   [25:0] id_router_022_src_channel;                                                                                      // id_router_022:src_channel -> rsp_xbar_demux_022:sink_channel
	wire          id_router_022_src_ready;                                                                                        // rsp_xbar_demux_022:sink_ready -> id_router_022:src_ready
	wire          cmd_xbar_demux_001_src23_ready;                                                                                 // PWM2_avalon_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src23_ready
	wire          id_router_023_src_endofpacket;                                                                                  // id_router_023:src_endofpacket -> rsp_xbar_demux_023:sink_endofpacket
	wire          id_router_023_src_valid;                                                                                        // id_router_023:src_valid -> rsp_xbar_demux_023:sink_valid
	wire          id_router_023_src_startofpacket;                                                                                // id_router_023:src_startofpacket -> rsp_xbar_demux_023:sink_startofpacket
	wire  [102:0] id_router_023_src_data;                                                                                         // id_router_023:src_data -> rsp_xbar_demux_023:sink_data
	wire   [25:0] id_router_023_src_channel;                                                                                      // id_router_023:src_channel -> rsp_xbar_demux_023:sink_channel
	wire          id_router_023_src_ready;                                                                                        // rsp_xbar_demux_023:sink_ready -> id_router_023:src_ready
	wire          cmd_xbar_demux_001_src24_ready;                                                                                 // PWM3_avalon_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src24_ready
	wire          id_router_024_src_endofpacket;                                                                                  // id_router_024:src_endofpacket -> rsp_xbar_demux_024:sink_endofpacket
	wire          id_router_024_src_valid;                                                                                        // id_router_024:src_valid -> rsp_xbar_demux_024:sink_valid
	wire          id_router_024_src_startofpacket;                                                                                // id_router_024:src_startofpacket -> rsp_xbar_demux_024:sink_startofpacket
	wire  [102:0] id_router_024_src_data;                                                                                         // id_router_024:src_data -> rsp_xbar_demux_024:sink_data
	wire   [25:0] id_router_024_src_channel;                                                                                      // id_router_024:src_channel -> rsp_xbar_demux_024:sink_channel
	wire          id_router_024_src_ready;                                                                                        // rsp_xbar_demux_024:sink_ready -> id_router_024:src_ready
	wire          cmd_xbar_demux_001_src25_ready;                                                                                 // pio_1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src25_ready
	wire          id_router_025_src_endofpacket;                                                                                  // id_router_025:src_endofpacket -> rsp_xbar_demux_025:sink_endofpacket
	wire          id_router_025_src_valid;                                                                                        // id_router_025:src_valid -> rsp_xbar_demux_025:sink_valid
	wire          id_router_025_src_startofpacket;                                                                                // id_router_025:src_startofpacket -> rsp_xbar_demux_025:sink_startofpacket
	wire  [102:0] id_router_025_src_data;                                                                                         // id_router_025:src_data -> rsp_xbar_demux_025:sink_data
	wire   [25:0] id_router_025_src_channel;                                                                                      // id_router_025:src_channel -> rsp_xbar_demux_025:sink_channel
	wire          id_router_025_src_ready;                                                                                        // rsp_xbar_demux_025:sink_ready -> id_router_025:src_ready
	wire          cmd_xbar_mux_001_src_endofpacket;                                                                               // cmd_xbar_mux_001:src_endofpacket -> width_adapter:in_endofpacket
	wire          cmd_xbar_mux_001_src_valid;                                                                                     // cmd_xbar_mux_001:src_valid -> width_adapter:in_valid
	wire          cmd_xbar_mux_001_src_startofpacket;                                                                             // cmd_xbar_mux_001:src_startofpacket -> width_adapter:in_startofpacket
	wire  [102:0] cmd_xbar_mux_001_src_data;                                                                                      // cmd_xbar_mux_001:src_data -> width_adapter:in_data
	wire   [25:0] cmd_xbar_mux_001_src_channel;                                                                                   // cmd_xbar_mux_001:src_channel -> width_adapter:in_channel
	wire          cmd_xbar_mux_001_src_ready;                                                                                     // width_adapter:in_ready -> cmd_xbar_mux_001:src_ready
	wire          width_adapter_src_endofpacket;                                                                                  // width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	wire          width_adapter_src_valid;                                                                                        // width_adapter:out_valid -> burst_adapter:sink0_valid
	wire          width_adapter_src_startofpacket;                                                                                // width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	wire   [84:0] width_adapter_src_data;                                                                                         // width_adapter:out_data -> burst_adapter:sink0_data
	wire          width_adapter_src_ready;                                                                                        // burst_adapter:sink0_ready -> width_adapter:out_ready
	wire   [25:0] width_adapter_src_channel;                                                                                      // width_adapter:out_channel -> burst_adapter:sink0_channel
	wire          id_router_001_src_endofpacket;                                                                                  // id_router_001:src_endofpacket -> width_adapter_001:in_endofpacket
	wire          id_router_001_src_valid;                                                                                        // id_router_001:src_valid -> width_adapter_001:in_valid
	wire          id_router_001_src_startofpacket;                                                                                // id_router_001:src_startofpacket -> width_adapter_001:in_startofpacket
	wire   [84:0] id_router_001_src_data;                                                                                         // id_router_001:src_data -> width_adapter_001:in_data
	wire   [25:0] id_router_001_src_channel;                                                                                      // id_router_001:src_channel -> width_adapter_001:in_channel
	wire          id_router_001_src_ready;                                                                                        // width_adapter_001:in_ready -> id_router_001:src_ready
	wire          width_adapter_001_src_endofpacket;                                                                              // width_adapter_001:out_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          width_adapter_001_src_valid;                                                                                    // width_adapter_001:out_valid -> rsp_xbar_demux_001:sink_valid
	wire          width_adapter_001_src_startofpacket;                                                                            // width_adapter_001:out_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [102:0] width_adapter_001_src_data;                                                                                     // width_adapter_001:out_data -> rsp_xbar_demux_001:sink_data
	wire          width_adapter_001_src_ready;                                                                                    // rsp_xbar_demux_001:sink_ready -> width_adapter_001:out_ready
	wire   [25:0] width_adapter_001_src_channel;                                                                                  // width_adapter_001:out_channel -> rsp_xbar_demux_001:sink_channel
	wire          crosser_out_endofpacket;                                                                                        // crosser:out_endofpacket -> adc_spi_read_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_out_valid;                                                                                              // crosser:out_valid -> adc_spi_read_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_out_startofpacket;                                                                                      // crosser:out_startofpacket -> adc_spi_read_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] crosser_out_data;                                                                                               // crosser:out_data -> adc_spi_read_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [25:0] crosser_out_channel;                                                                                            // crosser:out_channel -> adc_spi_read_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src11_endofpacket;                                                                           // cmd_xbar_demux_001:src11_endofpacket -> crosser:in_endofpacket
	wire          cmd_xbar_demux_001_src11_valid;                                                                                 // cmd_xbar_demux_001:src11_valid -> crosser:in_valid
	wire          cmd_xbar_demux_001_src11_startofpacket;                                                                         // cmd_xbar_demux_001:src11_startofpacket -> crosser:in_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src11_data;                                                                                  // cmd_xbar_demux_001:src11_data -> crosser:in_data
	wire   [25:0] cmd_xbar_demux_001_src11_channel;                                                                               // cmd_xbar_demux_001:src11_channel -> crosser:in_channel
	wire          cmd_xbar_demux_001_src11_ready;                                                                                 // crosser:in_ready -> cmd_xbar_demux_001:src11_ready
	wire          crosser_001_out_endofpacket;                                                                                    // crosser_001:out_endofpacket -> rsp_xbar_mux_001:sink11_endofpacket
	wire          crosser_001_out_valid;                                                                                          // crosser_001:out_valid -> rsp_xbar_mux_001:sink11_valid
	wire          crosser_001_out_startofpacket;                                                                                  // crosser_001:out_startofpacket -> rsp_xbar_mux_001:sink11_startofpacket
	wire  [102:0] crosser_001_out_data;                                                                                           // crosser_001:out_data -> rsp_xbar_mux_001:sink11_data
	wire   [25:0] crosser_001_out_channel;                                                                                        // crosser_001:out_channel -> rsp_xbar_mux_001:sink11_channel
	wire          crosser_001_out_ready;                                                                                          // rsp_xbar_mux_001:sink11_ready -> crosser_001:out_ready
	wire          rsp_xbar_demux_011_src0_endofpacket;                                                                            // rsp_xbar_demux_011:src0_endofpacket -> crosser_001:in_endofpacket
	wire          rsp_xbar_demux_011_src0_valid;                                                                                  // rsp_xbar_demux_011:src0_valid -> crosser_001:in_valid
	wire          rsp_xbar_demux_011_src0_startofpacket;                                                                          // rsp_xbar_demux_011:src0_startofpacket -> crosser_001:in_startofpacket
	wire  [102:0] rsp_xbar_demux_011_src0_data;                                                                                   // rsp_xbar_demux_011:src0_data -> crosser_001:in_data
	wire   [25:0] rsp_xbar_demux_011_src0_channel;                                                                                // rsp_xbar_demux_011:src0_channel -> crosser_001:in_channel
	wire          rsp_xbar_demux_011_src0_ready;                                                                                  // crosser_001:in_ready -> rsp_xbar_demux_011:src0_ready
	wire          irq_mapper_receiver0_irq;                                                                                       // timer:irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                                                                       // key:irq -> irq_mapper:receiver1_irq
	wire          irq_mapper_receiver2_irq;                                                                                       // sw:irq -> irq_mapper:receiver2_irq
	wire          irq_mapper_receiver3_irq;                                                                                       // jtag_uart_0:av_irq -> irq_mapper:receiver3_irq
	wire          irq_mapper_receiver4_irq;                                                                                       // uart_0:irq -> irq_mapper:receiver4_irq
	wire          irq_mapper_receiver5_irq;                                                                                       // epcs_flash_controller_0:irq -> irq_mapper:receiver5_irq
	wire   [31:0] nios2_qsys_0_d_irq_irq;                                                                                         // irq_mapper:sender_irq -> nios2_qsys_0:d_irq

	NIOS_Sys_nios2_qsys_0 nios2_qsys_0 (
		.clk                                   (altpll_0_c0_clk),                                                           //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                           //                   reset_n.reset_n
		.d_address                             (nios2_qsys_0_data_master_address),                                          //               data_master.address
		.d_byteenable                          (nios2_qsys_0_data_master_byteenable),                                       //                          .byteenable
		.d_read                                (nios2_qsys_0_data_master_read),                                             //                          .read
		.d_readdata                            (nios2_qsys_0_data_master_readdata),                                         //                          .readdata
		.d_waitrequest                         (nios2_qsys_0_data_master_waitrequest),                                      //                          .waitrequest
		.d_write                               (nios2_qsys_0_data_master_write),                                            //                          .write
		.d_writedata                           (nios2_qsys_0_data_master_writedata),                                        //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                                      //                          .debugaccess
		.i_address                             (nios2_qsys_0_instruction_master_address),                                   //        instruction_master.address
		.i_read                                (nios2_qsys_0_instruction_master_read),                                      //                          .read
		.i_readdata                            (nios2_qsys_0_instruction_master_readdata),                                  //                          .readdata
		.i_waitrequest                         (nios2_qsys_0_instruction_master_waitrequest),                               //                          .waitrequest
		.d_irq                                 (nios2_qsys_0_d_irq_irq),                                                    //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_0_jtag_debug_module_reset_reset),                                //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_read),        //                          .read
		.jtag_debug_module_readdata            (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write),       //                          .write
		.jtag_debug_module_writedata           (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                                           // custom_instruction_master.readra
	);

	NIOS_Sys_sdram sdram (
		.clk            (altpll_0_c0_clk),                                       //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),                   // reset.reset_n
		.az_addr        (sdram_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~sdram_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (sdram_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (sdram_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~sdram_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~sdram_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (sdram_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (sdram_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (sdram_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                                       //  wire.export
		.zs_ba          (sdram_wire_ba),                                         //      .export
		.zs_cas_n       (sdram_wire_cas_n),                                      //      .export
		.zs_cke         (sdram_wire_cke),                                        //      .export
		.zs_cs_n        (sdram_wire_cs_n),                                       //      .export
		.zs_dq          (sdram_wire_dq),                                         //      .export
		.zs_dqm         (sdram_wire_dqm),                                        //      .export
		.zs_ras_n       (sdram_wire_ras_n),                                      //      .export
		.zs_we_n        (sdram_wire_we_n)                                        //      .export
	);

	NIOS_Sys_led led (
		.clk        (altpll_0_c0_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),              //               reset.reset_n
		.address    (led_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~led_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (led_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (led_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (led_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (led_external_connection_export)                    // external_connection.export
	);

	NIOS_Sys_key key (
		.clk        (altpll_0_c0_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),              //               reset.reset_n
		.address    (key_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~key_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (key_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (key_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (key_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (key_external_connection_export),                   // external_connection.export
		.irq        (irq_mapper_receiver1_irq)                          //                 irq.irq
	);

	NIOS_Sys_sw sw (
		.clk        (altpll_0_c0_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),             //               reset.reset_n
		.address    (sw_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~sw_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (sw_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (sw_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (sw_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (sw_external_connection_export),                   // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                         //                 irq.irq
	);

	NIOS_Sys_timer timer (
		.clk        (altpll_0_c0_clk),                                    //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                // reset.reset_n
		.address    (timer_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                            //   irq.irq
	);

	NIOS_Sys_performance_counter performance_counter (
		.clk           (altpll_0_c0_clk),                                                                //           clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                                            //         reset.reset_n
		.address       (performance_counter_control_slave_translator_avalon_anti_slave_0_address),       // control_slave.address
		.begintransfer (performance_counter_control_slave_translator_avalon_anti_slave_0_begintransfer), //              .begintransfer
		.readdata      (performance_counter_control_slave_translator_avalon_anti_slave_0_readdata),      //              .readdata
		.write         (performance_counter_control_slave_translator_avalon_anti_slave_0_write),         //              .write
		.writedata     (performance_counter_control_slave_translator_avalon_anti_slave_0_writedata)      //              .writedata
	);

	NIOS_Sys_altpll_0 altpll_0 (
		.clk       (clk_clk),                            //       inclk_interface.clk
		.reset     (rst_controller_002_reset_out_reset), // inclk_interface_reset.reset
		.read      (),                                   //             pll_slave.read
		.write     (),                                   //                      .write
		.address   (),                                   //                      .address
		.readdata  (),                                   //                      .readdata
		.writedata (),                                   //                      .writedata
		.c0        (altpll_0_c0_clk),                    //                    c0.clk
		.c1        (altpll_0_c1_clk),                    //                    c1.clk
		.c2        (altpll_0_c2_clk),                    //                    c2.clk
		.areset    (),                                   //        areset_conduit.export
		.locked    (),                                   //        locked_conduit.export
		.phasedone ()                                    //     phasedone_conduit.export
	);

	Ultrasound_interface #(
		.idle             (5'b00001),
		.trigger          (5'b00010),
		.wait_feedback    (5'b00100),
		.measure_feedback (5'b01000)
	) ultrasound0 (
		.clk         (altpll_0_c0_clk),                                                      //          clock.clk
		.reset_n     (~rst_controller_001_reset_out_reset),                                  //          reset.reset_n
		.chipselect  (ultrasound0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), // avalon_slave_0.chipselect
		.address     (ultrasound0_avalon_slave_0_translator_avalon_anti_slave_0_address),    //               .address
		.write       (ultrasound0_avalon_slave_0_translator_avalon_anti_slave_0_write),      //               .write
		.writedata   (ultrasound0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),  //               .writedata
		.read        (ultrasound0_avalon_slave_0_translator_avalon_anti_slave_0_read),       //               .read
		.byteenable  (ultrasound0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable), //               .byteenable
		.readdata    (ultrasound0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),   //               .readdata
		.feedback_in (ultrasound0_conduit_end_feedback_in),                                  //    conduit_end.export
		.trigger_out (ultrasound0_conduit_end_trigger_out)                                   //               .export
	);

	Ultrasound_interface #(
		.idle             (5'b00001),
		.trigger          (5'b00010),
		.wait_feedback    (5'b00100),
		.measure_feedback (5'b01000)
	) ultrasound1 (
		.clk         (altpll_0_c0_clk),                                                      //          clock.clk
		.reset_n     (~rst_controller_001_reset_out_reset),                                  //          reset.reset_n
		.chipselect  (ultrasound1_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), // avalon_slave_0.chipselect
		.address     (ultrasound1_avalon_slave_0_translator_avalon_anti_slave_0_address),    //               .address
		.write       (ultrasound1_avalon_slave_0_translator_avalon_anti_slave_0_write),      //               .write
		.writedata   (ultrasound1_avalon_slave_0_translator_avalon_anti_slave_0_writedata),  //               .writedata
		.read        (ultrasound1_avalon_slave_0_translator_avalon_anti_slave_0_read),       //               .read
		.byteenable  (ultrasound1_avalon_slave_0_translator_avalon_anti_slave_0_byteenable), //               .byteenable
		.readdata    (ultrasound1_avalon_slave_0_translator_avalon_anti_slave_0_readdata),   //               .readdata
		.feedback_in (ultrasound1_conduit_end_feedback_in),                                  //    conduit_end.export
		.trigger_out (ultrasound1_conduit_end_trigger_out)                                   //               .export
	);

	TERASIC_ADC_READ adc_spi_read (
		.clk          (altpll_0_c2_clk),                                              //       clock.clk
		.reset_n      (~rst_controller_003_reset_out_reset),                          //       reset.reset_n
		.s_chipselect (adc_spi_read_slave_translator_avalon_anti_slave_0_chipselect), //       slave.chipselect
		.s_read       (adc_spi_read_slave_translator_avalon_anti_slave_0_read),       //            .read
		.s_readdata   (adc_spi_read_slave_translator_avalon_anti_slave_0_readdata),   //            .readdata
		.s_write      (adc_spi_read_slave_translator_avalon_anti_slave_0_write),      //            .write
		.s_writedata  (adc_spi_read_slave_translator_avalon_anti_slave_0_writedata),  //            .writedata
		.SPI_OUT      (adc_spi_read_conduit_end_OUT),                                 // conduit_end.export
		.SPI_IN       (adc_spi_read_conduit_end_IN),                                  //            .export
		.SPI_CS_n     (adc_spi_read_conduit_end_CS_n),                                //            .export
		.SPI_CLK      (adc_spi_read_conduit_end_CLK)                                  //            .export
	);

	pwm_gen pwm0 (
		.avs_address   (pwm0_avalon_slave_translator_avalon_anti_slave_0_address),    // avalon_slave.address
		.avs_write     (pwm0_avalon_slave_translator_avalon_anti_slave_0_write),      //             .write
		.avs_I_cs      (pwm0_avalon_slave_translator_avalon_anti_slave_0_chipselect), //             .chipselect
		.avs_I_wr_data (pwm0_avalon_slave_translator_avalon_anti_slave_0_writedata),  //             .writedata
		.csi_I_clk     (altpll_0_c0_clk),                                             //   clock_sink.clk
		.csi_I_rst     (~rst_controller_001_reset_out_reset),                         //  clock_reset.reset_n
		.coe_O_pwm1    (pwm0_conduit_end_pwm1),                                       //  conduit_end.export
		.coe_O_pwm2    (pwm0_conduit_end_pwm2)                                        //             .export
	);

	pwm_gen pwm1 (
		.avs_address   (pwm1_avalon_slave_translator_avalon_anti_slave_0_address),    // avalon_slave.address
		.avs_write     (pwm1_avalon_slave_translator_avalon_anti_slave_0_write),      //             .write
		.avs_I_cs      (pwm1_avalon_slave_translator_avalon_anti_slave_0_chipselect), //             .chipselect
		.avs_I_wr_data (pwm1_avalon_slave_translator_avalon_anti_slave_0_writedata),  //             .writedata
		.csi_I_clk     (altpll_0_c0_clk),                                             //   clock_sink.clk
		.csi_I_rst     (~rst_controller_001_reset_out_reset),                         //  clock_reset.reset_n
		.coe_O_pwm1    (pwm1_conduit_end_pwm1),                                       //  conduit_end.export
		.coe_O_pwm2    (pwm1_conduit_end_pwm2)                                        //             .export
	);

	NIOS_Sys_jtag_uart_0 jtag_uart_0 (
		.clk            (altpll_0_c0_clk),                                                          //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                                      //             reset.reset_n
		.av_chipselect  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver3_irq)                                                  //               irq.irq
	);

	pulse_senor_read encoder0 (
		.clk        (altpll_0_c0_clk),                                                   //          clock.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                               //          reset.reset_n
		.chipselect (encoder0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), // avalon_slave_0.chipselect
		.address    (encoder0_avalon_slave_0_translator_avalon_anti_slave_0_address),    //               .address
		.write      (encoder0_avalon_slave_0_translator_avalon_anti_slave_0_write),      //               .write
		.writedata  (encoder0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),  //               .writedata
		.read       (encoder0_avalon_slave_0_translator_avalon_anti_slave_0_read),       //               .read
		.readdata   (encoder0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),   //               .readdata
		.byteenable (encoder0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable), //               .byteenable
		.pulse_in   (encoder0_conduit_end_export)                                        //    conduit_end.export
	);

	pulse_senor_read encoder1 (
		.clk        (altpll_0_c0_clk),                                                   //          clock.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                               //          reset.reset_n
		.chipselect (encoder1_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), // avalon_slave_0.chipselect
		.address    (encoder1_avalon_slave_0_translator_avalon_anti_slave_0_address),    //               .address
		.write      (encoder1_avalon_slave_0_translator_avalon_anti_slave_0_write),      //               .write
		.writedata  (encoder1_avalon_slave_0_translator_avalon_anti_slave_0_writedata),  //               .writedata
		.read       (encoder1_avalon_slave_0_translator_avalon_anti_slave_0_read),       //               .read
		.readdata   (encoder1_avalon_slave_0_translator_avalon_anti_slave_0_readdata),   //               .readdata
		.byteenable (encoder1_avalon_slave_0_translator_avalon_anti_slave_0_byteenable), //               .byteenable
		.pulse_in   (encoder1_conduit_end_export)                                        //    conduit_end.export
	);

	NIOS_Sys_led pio_0 (
		.clk        (altpll_0_c0_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                //               reset.reset_n
		.address    (pio_0_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~pio_0_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (pio_0_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (pio_0_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (pio_0_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (pio_0_external_connection_export)                    // external_connection.export
	);

	NIOS_Sys_onchip_memory2_0 onchip_memory2_0 (
		.clk        (altpll_0_c0_clk),                                               //   clk1.clk
		.address    (onchip_memory2_0_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.clken      (onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.chipselect (onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.write      (onchip_memory2_0_s1_translator_avalon_anti_slave_0_write),      //       .write
		.readdata   (onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.writedata  (onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),                            // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req)                         //       .reset_req
	);

	NIOS_Sys_uart_0 uart_0 (
		.clk           (altpll_0_c0_clk),                                        //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                        //               reset.reset_n
		.address       (uart_0_s1_translator_avalon_anti_slave_0_address),       //                  s1.address
		.begintransfer (uart_0_s1_translator_avalon_anti_slave_0_begintransfer), //                    .begintransfer
		.chipselect    (uart_0_s1_translator_avalon_anti_slave_0_chipselect),    //                    .chipselect
		.read_n        (~uart_0_s1_translator_avalon_anti_slave_0_read),         //                    .read_n
		.write_n       (~uart_0_s1_translator_avalon_anti_slave_0_write),        //                    .write_n
		.writedata     (uart_0_s1_translator_avalon_anti_slave_0_writedata),     //                    .writedata
		.readdata      (uart_0_s1_translator_avalon_anti_slave_0_readdata),      //                    .readdata
		.dataavailable (),                                                       //                    .dataavailable
		.readyfordata  (),                                                       //                    .readyfordata
		.rxd           (uart_0_external_connection_rxd),                         // external_connection.export
		.txd           (uart_0_external_connection_txd),                         //                    .export
		.irq           (irq_mapper_receiver4_irq)                                //                 irq.irq
	);

	Ultrasound_interface #(
		.idle             (5'b00001),
		.trigger          (5'b00010),
		.wait_feedback    (5'b00100),
		.measure_feedback (5'b01000)
	) ultrasound2 (
		.clk         (altpll_0_c0_clk),                                                      //          clock.clk
		.reset_n     (~rst_controller_reset_out_reset),                                      //          reset.reset_n
		.chipselect  (ultrasound2_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), // avalon_slave_0.chipselect
		.address     (ultrasound2_avalon_slave_0_translator_avalon_anti_slave_0_address),    //               .address
		.write       (ultrasound2_avalon_slave_0_translator_avalon_anti_slave_0_write),      //               .write
		.writedata   (ultrasound2_avalon_slave_0_translator_avalon_anti_slave_0_writedata),  //               .writedata
		.read        (ultrasound2_avalon_slave_0_translator_avalon_anti_slave_0_read),       //               .read
		.byteenable  (ultrasound2_avalon_slave_0_translator_avalon_anti_slave_0_byteenable), //               .byteenable
		.readdata    (ultrasound2_avalon_slave_0_translator_avalon_anti_slave_0_readdata),   //               .readdata
		.feedback_in (ultrasound2_conduit_end_feedback_in),                                  //    conduit_end.export
		.trigger_out (ultrasound2_conduit_end_trigger_out)                                   //               .export
	);

	Ultrasound_interface #(
		.idle             (5'b00001),
		.trigger          (5'b00010),
		.wait_feedback    (5'b00100),
		.measure_feedback (5'b01000)
	) ultrasound3 (
		.clk         (altpll_0_c0_clk),                                                      //          clock.clk
		.reset_n     (~rst_controller_reset_out_reset),                                      //          reset.reset_n
		.chipselect  (ultrasound3_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), // avalon_slave_0.chipselect
		.address     (ultrasound3_avalon_slave_0_translator_avalon_anti_slave_0_address),    //               .address
		.write       (ultrasound3_avalon_slave_0_translator_avalon_anti_slave_0_write),      //               .write
		.writedata   (ultrasound3_avalon_slave_0_translator_avalon_anti_slave_0_writedata),  //               .writedata
		.read        (ultrasound3_avalon_slave_0_translator_avalon_anti_slave_0_read),       //               .read
		.byteenable  (ultrasound3_avalon_slave_0_translator_avalon_anti_slave_0_byteenable), //               .byteenable
		.readdata    (ultrasound3_avalon_slave_0_translator_avalon_anti_slave_0_readdata),   //               .readdata
		.feedback_in (ultrasound3_conduit_end_feedback_in),                                  //    conduit_end.export
		.trigger_out (ultrasound3_conduit_end_trigger_out)                                   //               .export
	);

	Ultrasound_interface #(
		.idle             (5'b00001),
		.trigger          (5'b00010),
		.wait_feedback    (5'b00100),
		.measure_feedback (5'b01000)
	) ultrasound4 (
		.clk         (altpll_0_c0_clk),                                                      //          clock.clk
		.reset_n     (~rst_controller_reset_out_reset),                                      //          reset.reset_n
		.chipselect  (ultrasound4_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), // avalon_slave_0.chipselect
		.address     (ultrasound4_avalon_slave_0_translator_avalon_anti_slave_0_address),    //               .address
		.write       (ultrasound4_avalon_slave_0_translator_avalon_anti_slave_0_write),      //               .write
		.writedata   (ultrasound4_avalon_slave_0_translator_avalon_anti_slave_0_writedata),  //               .writedata
		.read        (ultrasound4_avalon_slave_0_translator_avalon_anti_slave_0_read),       //               .read
		.byteenable  (ultrasound4_avalon_slave_0_translator_avalon_anti_slave_0_byteenable), //               .byteenable
		.readdata    (ultrasound4_avalon_slave_0_translator_avalon_anti_slave_0_readdata),   //               .readdata
		.feedback_in (ultrasound4_conduit_end_feedback_in),                                  //    conduit_end.export
		.trigger_out (ultrasound4_conduit_end_trigger_out)                                   //               .export
	);

	Ultrasound_interface #(
		.idle             (5'b00001),
		.trigger          (5'b00010),
		.wait_feedback    (5'b00100),
		.measure_feedback (5'b01000)
	) ultrasound5 (
		.clk         (altpll_0_c0_clk),                                                      //          clock.clk
		.reset_n     (~rst_controller_reset_out_reset),                                      //          reset.reset_n
		.chipselect  (ultrasound5_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), // avalon_slave_0.chipselect
		.address     (ultrasound5_avalon_slave_0_translator_avalon_anti_slave_0_address),    //               .address
		.write       (ultrasound5_avalon_slave_0_translator_avalon_anti_slave_0_write),      //               .write
		.writedata   (ultrasound5_avalon_slave_0_translator_avalon_anti_slave_0_writedata),  //               .writedata
		.read        (ultrasound5_avalon_slave_0_translator_avalon_anti_slave_0_read),       //               .read
		.byteenable  (ultrasound5_avalon_slave_0_translator_avalon_anti_slave_0_byteenable), //               .byteenable
		.readdata    (ultrasound5_avalon_slave_0_translator_avalon_anti_slave_0_readdata),   //               .readdata
		.feedback_in (ultrasound5_conduit_end_feedback_in),                                  //    conduit_end.export
		.trigger_out (ultrasound5_conduit_end_trigger_out)                                   //               .export
	);

	pwm_gen pwm2 (
		.avs_address   (pwm2_avalon_slave_translator_avalon_anti_slave_0_address),    // avalon_slave.address
		.avs_write     (pwm2_avalon_slave_translator_avalon_anti_slave_0_write),      //             .write
		.avs_I_cs      (pwm2_avalon_slave_translator_avalon_anti_slave_0_chipselect), //             .chipselect
		.avs_I_wr_data (pwm2_avalon_slave_translator_avalon_anti_slave_0_writedata),  //             .writedata
		.csi_I_clk     (altpll_0_c0_clk),                                             //   clock_sink.clk
		.csi_I_rst     (~rst_controller_reset_out_reset),                             //  clock_reset.reset_n
		.coe_O_pwm1    (pwm2_conduit_end_pwm1),                                       //  conduit_end.export
		.coe_O_pwm2    (pwm2_conduit_end_pwm2)                                        //             .export
	);

	pwm_gen pwm3 (
		.avs_address   (pwm3_avalon_slave_translator_avalon_anti_slave_0_address),    // avalon_slave.address
		.avs_write     (pwm3_avalon_slave_translator_avalon_anti_slave_0_write),      //             .write
		.avs_I_cs      (pwm3_avalon_slave_translator_avalon_anti_slave_0_chipselect), //             .chipselect
		.avs_I_wr_data (pwm3_avalon_slave_translator_avalon_anti_slave_0_writedata),  //             .writedata
		.csi_I_clk     (altpll_0_c0_clk),                                             //   clock_sink.clk
		.csi_I_rst     (~rst_controller_reset_out_reset),                             //  clock_reset.reset_n
		.coe_O_pwm1    (pwm3_conduit_end_pwm1),                                       //  conduit_end.export
		.coe_O_pwm2    (pwm3_conduit_end_pwm2)                                        //             .export
	);

	NIOS_Sys_pio_1 pio_1 (
		.clk      (altpll_0_c0_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address  (pio_1_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (pio_1_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (pio_1_external_connection_export)                  // external_connection.export
	);

	NIOS_Sys_epcs_flash_controller_0 epcs_flash_controller_0 (
		.clk           (altpll_0_c0_clk),                                                                     //               clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                                                     //             reset.reset_n
		.address       (epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_address),    // epcs_control_port.address
		.chipselect    (epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_chipselect), //                  .chipselect
		.dataavailable (),                                                                                    //                  .dataavailable
		.endofpacket   (),                                                                                    //                  .endofpacket
		.read_n        (~epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_read),      //                  .read_n
		.readdata      (epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_readdata),   //                  .readdata
		.readyfordata  (),                                                                                    //                  .readyfordata
		.write_n       (~epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_write),     //                  .write_n
		.writedata     (epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_writedata),  //                  .writedata
		.irq           (irq_mapper_receiver5_irq),                                                            //               irq.irq
		.dclk          (),                                                                                    //          external.export
		.sce           (),                                                                                    //                  .export
		.sdo           (),                                                                                    //                  .export
		.data0         ()                                                                                     //                  .export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (26),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (26),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_qsys_0_instruction_master_translator (
		.clk                      (altpll_0_c0_clk),                                                                    //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                     //                     reset.reset
		.uav_address              (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios2_qsys_0_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios2_qsys_0_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (nios2_qsys_0_instruction_master_read),                                               //                          .read
		.av_readdata              (nios2_qsys_0_instruction_master_readdata),                                           //                          .readdata
		.av_burstcount            (1'b1),                                                                               //               (terminated)
		.av_byteenable            (4'b1111),                                                                            //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                               //               (terminated)
		.av_begintransfer         (1'b0),                                                                               //               (terminated)
		.av_chipselect            (1'b0),                                                                               //               (terminated)
		.av_readdatavalid         (),                                                                                   //               (terminated)
		.av_write                 (1'b0),                                                                               //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                               //               (terminated)
		.av_lock                  (1'b0),                                                                               //               (terminated)
		.av_debugaccess           (1'b0),                                                                               //               (terminated)
		.uav_clken                (),                                                                                   //               (terminated)
		.av_clken                 (1'b1),                                                                               //               (terminated)
		.uav_response             (2'b00),                                                                              //               (terminated)
		.av_response              (),                                                                                   //               (terminated)
		.uav_writeresponserequest (),                                                                                   //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                               //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                               //               (terminated)
		.av_writeresponsevalid    ()                                                                                    //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (26),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (26),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (1)
	) nios2_qsys_0_data_master_translator (
		.clk                      (altpll_0_c0_clk),                                                             //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                              //                     reset.reset
		.uav_address              (nios2_qsys_0_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios2_qsys_0_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios2_qsys_0_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios2_qsys_0_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios2_qsys_0_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (nios2_qsys_0_data_master_byteenable),                                         //                          .byteenable
		.av_read                  (nios2_qsys_0_data_master_read),                                               //                          .read
		.av_readdata              (nios2_qsys_0_data_master_readdata),                                           //                          .readdata
		.av_write                 (nios2_qsys_0_data_master_write),                                              //                          .write
		.av_writedata             (nios2_qsys_0_data_master_writedata),                                          //                          .writedata
		.av_debugaccess           (nios2_qsys_0_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount            (1'b1),                                                                        //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                        //               (terminated)
		.av_begintransfer         (1'b0),                                                                        //               (terminated)
		.av_chipselect            (1'b0),                                                                        //               (terminated)
		.av_readdatavalid         (),                                                                            //               (terminated)
		.av_lock                  (1'b0),                                                                        //               (terminated)
		.uav_clken                (),                                                                            //               (terminated)
		.av_clken                 (1'b1),                                                                        //               (terminated)
		.uav_response             (2'b00),                                                                       //               (terminated)
		.av_response              (),                                                                            //               (terminated)
		.uav_writeresponserequest (),                                                                            //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                        //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                        //               (terminated)
		.av_writeresponsevalid    ()                                                                             //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) nios2_qsys_0_jtag_debug_module_translator (
		.clk                      (altpll_0_c0_clk),                                                                           //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                            //                    reset.reset
		.uav_address              (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                                          //              (terminated)
		.av_burstcount            (),                                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                                          //              (terminated)
		.av_lock                  (),                                                                                          //              (terminated)
		.av_chipselect            (),                                                                                          //              (terminated)
		.av_clken                 (),                                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                                      //              (terminated)
		.av_outputenable          (),                                                                                          //              (terminated)
		.uav_response             (),                                                                                          //              (terminated)
		.av_response              (2'b00),                                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (24),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sdram_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                     //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                  //                    reset.reset
		.uav_address              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sdram_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (sdram_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (sdram_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (sdram_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (sdram_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (sdram_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (sdram_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (sdram_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (sdram_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (12),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_memory2_0_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                                //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                             //                    reset.reset
		.uav_address              (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (onchip_memory2_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (onchip_memory2_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken                 (onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read                  (),                                                                               //              (terminated)
		.av_begintransfer         (),                                                                               //              (terminated)
		.av_beginbursttransfer    (),                                                                               //              (terminated)
		.av_burstcount            (),                                                                               //              (terminated)
		.av_readdatavalid         (1'b0),                                                                           //              (terminated)
		.av_waitrequest           (1'b0),                                                                           //              (terminated)
		.av_writebyteenable       (),                                                                               //              (terminated)
		.av_lock                  (),                                                                               //              (terminated)
		.uav_clken                (1'b0),                                                                           //              (terminated)
		.av_debugaccess           (),                                                                               //              (terminated)
		.av_outputenable          (),                                                                               //              (terminated)
		.uav_response             (),                                                                               //              (terminated)
		.av_response              (2'b00),                                                                          //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                           //              (terminated)
		.uav_writeresponsevalid   (),                                                                               //              (terminated)
		.av_writeresponserequest  (),                                                                               //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) epcs_flash_controller_0_epcs_control_port_translator (
		.clk                      (altpll_0_c0_clk),                                                                                      //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                                       //                    reset.reset
		.uav_address              (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                                     //              (terminated)
		.av_beginbursttransfer    (),                                                                                                     //              (terminated)
		.av_burstcount            (),                                                                                                     //              (terminated)
		.av_byteenable            (),                                                                                                     //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                                 //              (terminated)
		.av_waitrequest           (1'b0),                                                                                                 //              (terminated)
		.av_writebyteenable       (),                                                                                                     //              (terminated)
		.av_lock                  (),                                                                                                     //              (terminated)
		.av_clken                 (),                                                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                                                 //              (terminated)
		.av_debugaccess           (),                                                                                                     //              (terminated)
		.av_outputenable          (),                                                                                                     //              (terminated)
		.uav_response             (),                                                                                                     //              (terminated)
		.av_response              (2'b00),                                                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) led_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                   //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                //                    reset.reset
		.uav_address              (led_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (led_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (led_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (led_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (led_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (led_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (led_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (led_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (led_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (led_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (led_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                  //              (terminated)
		.av_begintransfer         (),                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                  //              (terminated)
		.av_burstcount            (),                                                                  //              (terminated)
		.av_byteenable            (),                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                              //              (terminated)
		.av_waitrequest           (1'b0),                                                              //              (terminated)
		.av_writebyteenable       (),                                                                  //              (terminated)
		.av_lock                  (),                                                                  //              (terminated)
		.av_clken                 (),                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                              //              (terminated)
		.av_debugaccess           (),                                                                  //              (terminated)
		.av_outputenable          (),                                                                  //              (terminated)
		.uav_response             (),                                                                  //              (terminated)
		.av_response              (2'b00),                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) key_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                   //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                //                    reset.reset
		.uav_address              (key_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (key_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (key_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (key_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (key_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (key_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (key_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (key_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (key_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (key_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (key_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (key_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (key_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (key_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (key_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (key_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                  //              (terminated)
		.av_begintransfer         (),                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                  //              (terminated)
		.av_burstcount            (),                                                                  //              (terminated)
		.av_byteenable            (),                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                              //              (terminated)
		.av_waitrequest           (1'b0),                                                              //              (terminated)
		.av_writebyteenable       (),                                                                  //              (terminated)
		.av_lock                  (),                                                                  //              (terminated)
		.av_clken                 (),                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                              //              (terminated)
		.av_debugaccess           (),                                                                  //              (terminated)
		.av_outputenable          (),                                                                  //              (terminated)
		.uav_response             (),                                                                  //              (terminated)
		.av_response              (2'b00),                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sw_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                               //                    reset.reset
		.uav_address              (sw_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sw_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sw_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sw_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sw_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sw_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sw_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (sw_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (sw_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (sw_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (sw_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                 //              (terminated)
		.av_begintransfer         (),                                                                 //              (terminated)
		.av_beginbursttransfer    (),                                                                 //              (terminated)
		.av_burstcount            (),                                                                 //              (terminated)
		.av_byteenable            (),                                                                 //              (terminated)
		.av_readdatavalid         (1'b0),                                                             //              (terminated)
		.av_waitrequest           (1'b0),                                                             //              (terminated)
		.av_writebyteenable       (),                                                                 //              (terminated)
		.av_lock                  (),                                                                 //              (terminated)
		.av_clken                 (),                                                                 //              (terminated)
		.uav_clken                (1'b0),                                                             //              (terminated)
		.av_debugaccess           (),                                                                 //              (terminated)
		.av_outputenable          (),                                                                 //              (terminated)
		.uav_response             (),                                                                 //              (terminated)
		.av_response              (2'b00),                                                            //              (terminated)
		.uav_writeresponserequest (1'b0),                                                             //              (terminated)
		.uav_writeresponsevalid   (),                                                                 //              (terminated)
		.av_writeresponserequest  (),                                                                 //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                     //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                  //                    reset.reset
		.uav_address              (timer_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (timer_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (timer_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (timer_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (timer_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (timer_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (timer_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                    //              (terminated)
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_byteenable            (),                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (4),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) performance_counter_control_slave_translator (
		.clk                      (altpll_0_c0_clk),                                                                              //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                           //                    reset.reset
		.uav_address              (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (performance_counter_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (performance_counter_control_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (performance_counter_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (performance_counter_control_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (performance_counter_control_slave_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_read                  (),                                                                                             //              (terminated)
		.av_beginbursttransfer    (),                                                                                             //              (terminated)
		.av_burstcount            (),                                                                                             //              (terminated)
		.av_byteenable            (),                                                                                             //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                         //              (terminated)
		.av_waitrequest           (1'b0),                                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                                             //              (terminated)
		.av_lock                  (),                                                                                             //              (terminated)
		.av_chipselect            (),                                                                                             //              (terminated)
		.av_clken                 (),                                                                                             //              (terminated)
		.uav_clken                (1'b0),                                                                                         //              (terminated)
		.av_debugaccess           (),                                                                                             //              (terminated)
		.av_outputenable          (),                                                                                             //              (terminated)
		.uav_response             (),                                                                                             //              (terminated)
		.av_response              (2'b00),                                                                                        //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                         //              (terminated)
		.uav_writeresponsevalid   (),                                                                                             //              (terminated)
		.av_writeresponserequest  (),                                                                                             //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ultrasound0_avalon_slave_0_translator (
		.clk                      (altpll_0_c0_clk),                                                                       //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                    //                    reset.reset
		.uav_address              (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ultrasound0_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ultrasound0_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (ultrasound0_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (ultrasound0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ultrasound0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (ultrasound0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (ultrasound0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                                      //              (terminated)
		.av_burstcount            (),                                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                                      //              (terminated)
		.av_lock                  (),                                                                                      //              (terminated)
		.av_clken                 (),                                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                                  //              (terminated)
		.av_debugaccess           (),                                                                                      //              (terminated)
		.av_outputenable          (),                                                                                      //              (terminated)
		.uav_response             (),                                                                                      //              (terminated)
		.av_response              (2'b00),                                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ultrasound1_avalon_slave_0_translator (
		.clk                      (altpll_0_c0_clk),                                                                       //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                    //                    reset.reset
		.uav_address              (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ultrasound1_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ultrasound1_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (ultrasound1_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (ultrasound1_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ultrasound1_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (ultrasound1_avalon_slave_0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (ultrasound1_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                                      //              (terminated)
		.av_burstcount            (),                                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                                      //              (terminated)
		.av_lock                  (),                                                                                      //              (terminated)
		.av_clken                 (),                                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                                  //              (terminated)
		.av_debugaccess           (),                                                                                      //              (terminated)
		.av_outputenable          (),                                                                                      //              (terminated)
		.uav_response             (),                                                                                      //              (terminated)
		.av_response              (2'b00),                                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) adc_spi_read_slave_translator (
		.clk                      (altpll_0_c2_clk),                                                               //                      clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                            //                    reset.reset
		.uav_address              (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write                 (adc_spi_read_slave_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read                  (adc_spi_read_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (adc_spi_read_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (adc_spi_read_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (adc_spi_read_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_address               (),                                                                              //              (terminated)
		.av_begintransfer         (),                                                                              //              (terminated)
		.av_beginbursttransfer    (),                                                                              //              (terminated)
		.av_burstcount            (),                                                                              //              (terminated)
		.av_byteenable            (),                                                                              //              (terminated)
		.av_readdatavalid         (1'b0),                                                                          //              (terminated)
		.av_waitrequest           (1'b0),                                                                          //              (terminated)
		.av_writebyteenable       (),                                                                              //              (terminated)
		.av_lock                  (),                                                                              //              (terminated)
		.av_clken                 (),                                                                              //              (terminated)
		.uav_clken                (1'b0),                                                                          //              (terminated)
		.av_debugaccess           (),                                                                              //              (terminated)
		.av_outputenable          (),                                                                              //              (terminated)
		.uav_response             (),                                                                              //              (terminated)
		.av_response              (2'b00),                                                                         //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                          //              (terminated)
		.uav_writeresponsevalid   (),                                                                              //              (terminated)
		.av_writeresponserequest  (),                                                                              //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pwm0_avalon_slave_translator (
		.clk                      (altpll_0_c0_clk),                                                              //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                           //                    reset.reset
		.uav_address              (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (pwm0_avalon_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (pwm0_avalon_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_writedata             (pwm0_avalon_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (pwm0_avalon_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                             //              (terminated)
		.av_readdata              (32'b11011110101011011101111010101101),                                         //              (terminated)
		.av_begintransfer         (),                                                                             //              (terminated)
		.av_beginbursttransfer    (),                                                                             //              (terminated)
		.av_burstcount            (),                                                                             //              (terminated)
		.av_byteenable            (),                                                                             //              (terminated)
		.av_readdatavalid         (1'b0),                                                                         //              (terminated)
		.av_waitrequest           (1'b0),                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                             //              (terminated)
		.av_lock                  (),                                                                             //              (terminated)
		.av_clken                 (),                                                                             //              (terminated)
		.uav_clken                (1'b0),                                                                         //              (terminated)
		.av_debugaccess           (),                                                                             //              (terminated)
		.av_outputenable          (),                                                                             //              (terminated)
		.uav_response             (),                                                                             //              (terminated)
		.av_response              (2'b00),                                                                        //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                         //              (terminated)
		.uav_writeresponsevalid   (),                                                                             //              (terminated)
		.av_writeresponserequest  (),                                                                             //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pwm1_avalon_slave_translator (
		.clk                      (altpll_0_c0_clk),                                                              //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                           //                    reset.reset
		.uav_address              (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (pwm1_avalon_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (pwm1_avalon_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_writedata             (pwm1_avalon_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (pwm1_avalon_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                             //              (terminated)
		.av_readdata              (32'b11011110101011011101111010101101),                                         //              (terminated)
		.av_begintransfer         (),                                                                             //              (terminated)
		.av_beginbursttransfer    (),                                                                             //              (terminated)
		.av_burstcount            (),                                                                             //              (terminated)
		.av_byteenable            (),                                                                             //              (terminated)
		.av_readdatavalid         (1'b0),                                                                         //              (terminated)
		.av_waitrequest           (1'b0),                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                             //              (terminated)
		.av_lock                  (),                                                                             //              (terminated)
		.av_clken                 (),                                                                             //              (terminated)
		.uav_clken                (1'b0),                                                                         //              (terminated)
		.av_debugaccess           (),                                                                             //              (terminated)
		.av_outputenable          (),                                                                             //              (terminated)
		.uav_response             (),                                                                             //              (terminated)
		.av_response              (2'b00),                                                                        //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                         //              (terminated)
		.uav_writeresponsevalid   (),                                                                             //              (terminated)
		.av_writeresponserequest  (),                                                                             //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_0_avalon_jtag_slave_translator (
		.clk                      (altpll_0_c0_clk),                                                                          //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                       //                    reset.reset
		.uav_address              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                                         //              (terminated)
		.av_burstcount            (),                                                                                         //              (terminated)
		.av_byteenable            (),                                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                                         //              (terminated)
		.av_lock                  (),                                                                                         //              (terminated)
		.av_clken                 (),                                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                                     //              (terminated)
		.av_debugaccess           (),                                                                                         //              (terminated)
		.av_outputenable          (),                                                                                         //              (terminated)
		.uav_response             (),                                                                                         //              (terminated)
		.av_response              (2'b00),                                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (2),
		.AV_WRITE_WAIT_CYCLES           (2),
		.AV_SETUP_WAIT_CYCLES           (1),
		.AV_DATA_HOLD_CYCLES            (2)
	) encoder0_avalon_slave_0_translator (
		.clk                      (altpll_0_c0_clk),                                                                    //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                 //                    reset.reset
		.uav_address              (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (encoder0_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (encoder0_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (encoder0_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (encoder0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (encoder0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (encoder0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (encoder0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                                   //              (terminated)
		.av_burstcount            (),                                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                                               //              (terminated)
		.av_writebyteenable       (),                                                                                   //              (terminated)
		.av_lock                  (),                                                                                   //              (terminated)
		.av_clken                 (),                                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                                               //              (terminated)
		.av_debugaccess           (),                                                                                   //              (terminated)
		.av_outputenable          (),                                                                                   //              (terminated)
		.uav_response             (),                                                                                   //              (terminated)
		.av_response              (2'b00),                                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (2),
		.AV_WRITE_WAIT_CYCLES           (2),
		.AV_SETUP_WAIT_CYCLES           (1),
		.AV_DATA_HOLD_CYCLES            (2)
	) encoder1_avalon_slave_0_translator (
		.clk                      (altpll_0_c0_clk),                                                                    //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                 //                    reset.reset
		.uav_address              (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (encoder1_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (encoder1_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (encoder1_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (encoder1_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (encoder1_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (encoder1_avalon_slave_0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (encoder1_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                                   //              (terminated)
		.av_burstcount            (),                                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                                               //              (terminated)
		.av_writebyteenable       (),                                                                                   //              (terminated)
		.av_lock                  (),                                                                                   //              (terminated)
		.av_clken                 (),                                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                                               //              (terminated)
		.av_debugaccess           (),                                                                                   //              (terminated)
		.av_outputenable          (),                                                                                   //              (terminated)
		.uav_response             (),                                                                                   //              (terminated)
		.av_response              (2'b00),                                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pio_0_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                     //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                  //                    reset.reset
		.uav_address              (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (pio_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (pio_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (pio_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (pio_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (pio_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                    //              (terminated)
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_byteenable            (),                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) uart_0_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                      //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                       //                    reset.reset
		.uav_address              (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (uart_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (uart_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (uart_0_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (uart_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (uart_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (uart_0_s1_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_chipselect            (uart_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_beginbursttransfer    (),                                                                     //              (terminated)
		.av_burstcount            (),                                                                     //              (terminated)
		.av_byteenable            (),                                                                     //              (terminated)
		.av_readdatavalid         (1'b0),                                                                 //              (terminated)
		.av_waitrequest           (1'b0),                                                                 //              (terminated)
		.av_writebyteenable       (),                                                                     //              (terminated)
		.av_lock                  (),                                                                     //              (terminated)
		.av_clken                 (),                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                 //              (terminated)
		.av_debugaccess           (),                                                                     //              (terminated)
		.av_outputenable          (),                                                                     //              (terminated)
		.uav_response             (),                                                                     //              (terminated)
		.av_response              (2'b00),                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ultrasound2_avalon_slave_0_translator (
		.clk                      (altpll_0_c0_clk),                                                                       //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                        //                    reset.reset
		.uav_address              (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ultrasound2_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ultrasound2_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (ultrasound2_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (ultrasound2_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ultrasound2_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (ultrasound2_avalon_slave_0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (ultrasound2_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                                      //              (terminated)
		.av_burstcount            (),                                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                                      //              (terminated)
		.av_lock                  (),                                                                                      //              (terminated)
		.av_clken                 (),                                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                                  //              (terminated)
		.av_debugaccess           (),                                                                                      //              (terminated)
		.av_outputenable          (),                                                                                      //              (terminated)
		.uav_response             (),                                                                                      //              (terminated)
		.av_response              (2'b00),                                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ultrasound3_avalon_slave_0_translator (
		.clk                      (altpll_0_c0_clk),                                                                       //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                        //                    reset.reset
		.uav_address              (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ultrasound3_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ultrasound3_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (ultrasound3_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (ultrasound3_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ultrasound3_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (ultrasound3_avalon_slave_0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (ultrasound3_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                                      //              (terminated)
		.av_burstcount            (),                                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                                      //              (terminated)
		.av_lock                  (),                                                                                      //              (terminated)
		.av_clken                 (),                                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                                  //              (terminated)
		.av_debugaccess           (),                                                                                      //              (terminated)
		.av_outputenable          (),                                                                                      //              (terminated)
		.uav_response             (),                                                                                      //              (terminated)
		.av_response              (2'b00),                                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ultrasound4_avalon_slave_0_translator (
		.clk                      (altpll_0_c0_clk),                                                                       //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                        //                    reset.reset
		.uav_address              (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ultrasound4_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ultrasound4_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (ultrasound4_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (ultrasound4_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ultrasound4_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (ultrasound4_avalon_slave_0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (ultrasound4_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                                      //              (terminated)
		.av_burstcount            (),                                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                                      //              (terminated)
		.av_lock                  (),                                                                                      //              (terminated)
		.av_clken                 (),                                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                                  //              (terminated)
		.av_debugaccess           (),                                                                                      //              (terminated)
		.av_outputenable          (),                                                                                      //              (terminated)
		.uav_response             (),                                                                                      //              (terminated)
		.av_response              (2'b00),                                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ultrasound5_avalon_slave_0_translator (
		.clk                      (altpll_0_c0_clk),                                                                       //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                        //                    reset.reset
		.uav_address              (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ultrasound5_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ultrasound5_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (ultrasound5_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (ultrasound5_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ultrasound5_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (ultrasound5_avalon_slave_0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (ultrasound5_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                                      //              (terminated)
		.av_burstcount            (),                                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                                      //              (terminated)
		.av_lock                  (),                                                                                      //              (terminated)
		.av_clken                 (),                                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                                  //              (terminated)
		.av_debugaccess           (),                                                                                      //              (terminated)
		.av_outputenable          (),                                                                                      //              (terminated)
		.uav_response             (),                                                                                      //              (terminated)
		.av_response              (2'b00),                                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pwm2_avalon_slave_translator (
		.clk                      (altpll_0_c0_clk),                                                              //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                               //                    reset.reset
		.uav_address              (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (pwm2_avalon_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (pwm2_avalon_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_writedata             (pwm2_avalon_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (pwm2_avalon_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                             //              (terminated)
		.av_readdata              (32'b11011110101011011101111010101101),                                         //              (terminated)
		.av_begintransfer         (),                                                                             //              (terminated)
		.av_beginbursttransfer    (),                                                                             //              (terminated)
		.av_burstcount            (),                                                                             //              (terminated)
		.av_byteenable            (),                                                                             //              (terminated)
		.av_readdatavalid         (1'b0),                                                                         //              (terminated)
		.av_waitrequest           (1'b0),                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                             //              (terminated)
		.av_lock                  (),                                                                             //              (terminated)
		.av_clken                 (),                                                                             //              (terminated)
		.uav_clken                (1'b0),                                                                         //              (terminated)
		.av_debugaccess           (),                                                                             //              (terminated)
		.av_outputenable          (),                                                                             //              (terminated)
		.uav_response             (),                                                                             //              (terminated)
		.av_response              (2'b00),                                                                        //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                         //              (terminated)
		.uav_writeresponsevalid   (),                                                                             //              (terminated)
		.av_writeresponserequest  (),                                                                             //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pwm3_avalon_slave_translator (
		.clk                      (altpll_0_c0_clk),                                                              //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                               //                    reset.reset
		.uav_address              (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (pwm3_avalon_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (pwm3_avalon_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_writedata             (pwm3_avalon_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (pwm3_avalon_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                             //              (terminated)
		.av_readdata              (32'b11011110101011011101111010101101),                                         //              (terminated)
		.av_begintransfer         (),                                                                             //              (terminated)
		.av_beginbursttransfer    (),                                                                             //              (terminated)
		.av_burstcount            (),                                                                             //              (terminated)
		.av_byteenable            (),                                                                             //              (terminated)
		.av_readdatavalid         (1'b0),                                                                         //              (terminated)
		.av_waitrequest           (1'b0),                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                             //              (terminated)
		.av_lock                  (),                                                                             //              (terminated)
		.av_clken                 (),                                                                             //              (terminated)
		.uav_clken                (1'b0),                                                                         //              (terminated)
		.av_debugaccess           (),                                                                             //              (terminated)
		.av_outputenable          (),                                                                             //              (terminated)
		.uav_response             (),                                                                             //              (terminated)
		.av_response              (2'b00),                                                                        //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                         //              (terminated)
		.uav_writeresponsevalid   (),                                                                             //              (terminated)
		.av_writeresponserequest  (),                                                                             //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pio_1_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                     //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                      //                    reset.reset
		.uav_address              (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (pio_1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (pio_1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                    //              (terminated)
		.av_read                  (),                                                                    //              (terminated)
		.av_writedata             (),                                                                    //              (terminated)
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_byteenable            (),                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_chipselect            (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_BEGIN_BURST           (81),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.PKT_BURST_TYPE_H          (78),
		.PKT_BURST_TYPE_L          (77),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_TRANS_EXCLUSIVE       (67),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_THREAD_ID_H           (93),
		.PKT_THREAD_ID_L           (93),
		.PKT_CACHE_H               (100),
		.PKT_CACHE_L               (97),
		.PKT_DATA_SIDEBAND_H       (80),
		.PKT_DATA_SIDEBAND_L       (80),
		.PKT_QOS_H                 (82),
		.PKT_QOS_L                 (82),
		.PKT_ADDR_SIDEBAND_H       (79),
		.PKT_ADDR_SIDEBAND_L       (79),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.ST_DATA_W                 (103),
		.ST_CHANNEL_W              (26),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                             //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.av_address              (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_src_valid),                                                                      //        rp.valid
		.rp_data                 (rsp_xbar_mux_src_data),                                                                       //          .data
		.rp_channel              (rsp_xbar_mux_src_channel),                                                                    //          .channel
		.rp_startofpacket        (rsp_xbar_mux_src_startofpacket),                                                              //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_src_endofpacket),                                                                //          .endofpacket
		.rp_ready                (rsp_xbar_mux_src_ready),                                                                      //          .ready
		.av_response             (),                                                                                            // (terminated)
		.av_writeresponserequest (1'b0),                                                                                        // (terminated)
		.av_writeresponsevalid   ()                                                                                             // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_BEGIN_BURST           (81),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.PKT_BURST_TYPE_H          (78),
		.PKT_BURST_TYPE_L          (77),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_TRANS_EXCLUSIVE       (67),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_THREAD_ID_H           (93),
		.PKT_THREAD_ID_L           (93),
		.PKT_CACHE_H               (100),
		.PKT_CACHE_L               (97),
		.PKT_DATA_SIDEBAND_H       (80),
		.PKT_DATA_SIDEBAND_L       (80),
		.PKT_QOS_H                 (82),
		.PKT_QOS_L                 (82),
		.PKT_ADDR_SIDEBAND_H       (79),
		.PKT_ADDR_SIDEBAND_L       (79),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.ST_DATA_W                 (103),
		.ST_CHANNEL_W              (26),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                      //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.av_address              (nios2_qsys_0_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios2_qsys_0_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios2_qsys_0_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_001_src_valid),                                                           //        rp.valid
		.rp_data                 (rsp_xbar_mux_001_src_data),                                                            //          .data
		.rp_channel              (rsp_xbar_mux_001_src_channel),                                                         //          .channel
		.rp_startofpacket        (rsp_xbar_mux_001_src_startofpacket),                                                   //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_001_src_endofpacket),                                                     //          .endofpacket
		.rp_ready                (rsp_xbar_mux_001_src_ready),                                                           //          .ready
		.av_response             (),                                                                                     // (terminated)
		.av_writeresponserequest (1'b0),                                                                                 // (terminated)
		.av_writeresponsevalid   ()                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                                     //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                      //       clk_reset.reset
		.m0_address              (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                              //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                              //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                               //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                            //                .channel
		.rf_sink_ready           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                      // clk_reset.reset
		.in_data           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                                // (terminated)
		.csr_readdata      (),                                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                // (terminated)
		.almost_full_data  (),                                                                                                    // (terminated)
		.almost_empty_data (),                                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                                // (terminated)
		.out_empty         (),                                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                                // (terminated)
		.out_error         (),                                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                                // (terminated)
		.out_channel       ()                                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (43),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (44),
		.PKT_TRANS_POSTED          (45),
		.PKT_TRANS_WRITE           (46),
		.PKT_TRANS_READ            (47),
		.PKT_TRANS_LOCK            (48),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (53),
		.PKT_BYTE_CNT_H            (52),
		.PKT_BYTE_CNT_L            (50),
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (85),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                               //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                            //       clk_reset.reset
		.m0_address              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                   //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                   //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                    //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                             //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                 //                .channel
		.rf_sink_ready           (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (86),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                               //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.in_data           (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (18),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c0_clk),                                                         //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.in_data           (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                   // (terminated)
		.csr_read          (1'b0),                                                                    // (terminated)
		.csr_write         (1'b0),                                                                    // (terminated)
		.csr_readdata      (),                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                    // (terminated)
		.almost_full_data  (),                                                                        // (terminated)
		.almost_empty_data (),                                                                        // (terminated)
		.in_startofpacket  (1'b0),                                                                    // (terminated)
		.in_endofpacket    (1'b0),                                                                    // (terminated)
		.out_startofpacket (),                                                                        // (terminated)
		.out_endofpacket   (),                                                                        // (terminated)
		.in_empty          (1'b0),                                                                    // (terminated)
		.out_empty         (),                                                                        // (terminated)
		.in_error          (1'b0),                                                                    // (terminated)
		.out_error         (),                                                                        // (terminated)
		.in_channel        (1'b0),                                                                    // (terminated)
		.out_channel       ()                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_002_src_ready),                                                               //              cp.ready
		.cp_valid                (cmd_xbar_mux_002_src_valid),                                                               //                .valid
		.cp_data                 (cmd_xbar_mux_002_src_data),                                                                //                .data
		.cp_startofpacket        (cmd_xbar_mux_002_src_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_002_src_endofpacket),                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_mux_002_src_channel),                                                             //                .channel
		.rf_sink_ready           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                    //     (terminated)
		.m0_writeresponserequest (),                                                                                         //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                      //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                          //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                                 //       clk_reset.reset
		.m0_address              (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_003_src_ready),                                                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_003_src_valid),                                                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_003_src_data),                                                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_003_src_startofpacket),                                                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_003_src_endofpacket),                                                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_003_src_channel),                                                                                   //                .channel
		.rf_sink_ready           (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                                 // clk_reset.reset
		.in_data           (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                          // (terminated)
		.csr_read          (1'b0),                                                                                                           // (terminated)
		.csr_write         (1'b0),                                                                                                           // (terminated)
		.csr_readdata      (),                                                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                           // (terminated)
		.almost_full_data  (),                                                                                                               // (terminated)
		.almost_empty_data (),                                                                                                               // (terminated)
		.in_empty          (1'b0),                                                                                                           // (terminated)
		.out_empty         (),                                                                                                               // (terminated)
		.in_error          (1'b0),                                                                                                           // (terminated)
		.out_error         (),                                                                                                               // (terminated)
		.in_channel        (1'b0),                                                                                                           // (terminated)
		.out_channel       ()                                                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) led_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                          //       clk_reset.reset
		.m0_address              (led_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (led_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (led_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (led_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (led_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (led_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (led_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (led_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (led_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src4_ready),                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src4_valid),                                               //                .valid
		.cp_data                 (cmd_xbar_demux_001_src4_data),                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src4_startofpacket),                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src4_endofpacket),                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src4_channel),                                             //                .channel
		.rf_sink_ready           (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (led_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.in_data           (led_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                       // (terminated)
		.csr_read          (1'b0),                                                                        // (terminated)
		.csr_write         (1'b0),                                                                        // (terminated)
		.csr_readdata      (),                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                        // (terminated)
		.almost_full_data  (),                                                                            // (terminated)
		.almost_empty_data (),                                                                            // (terminated)
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_channel        (1'b0),                                                                        // (terminated)
		.out_channel       ()                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) key_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                          //       clk_reset.reset
		.m0_address              (key_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (key_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (key_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (key_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (key_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (key_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (key_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (key_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (key_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (key_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (key_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (key_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (key_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (key_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (key_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (key_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src5_ready),                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src5_valid),                                               //                .valid
		.cp_data                 (cmd_xbar_demux_001_src5_data),                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src5_startofpacket),                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src5_endofpacket),                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src5_channel),                                             //                .channel
		.rf_sink_ready           (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (key_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (key_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (key_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (key_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (key_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.in_data           (key_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (key_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (key_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (key_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (key_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                       // (terminated)
		.csr_read          (1'b0),                                                                        // (terminated)
		.csr_write         (1'b0),                                                                        // (terminated)
		.csr_readdata      (),                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                        // (terminated)
		.almost_full_data  (),                                                                            // (terminated)
		.almost_empty_data (),                                                                            // (terminated)
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_channel        (1'b0),                                                                        // (terminated)
		.out_channel       ()                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sw_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                         //       clk_reset.reset
		.m0_address              (sw_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sw_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sw_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sw_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sw_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sw_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sw_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sw_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sw_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src6_ready),                                              //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src6_valid),                                              //                .valid
		.cp_data                 (cmd_xbar_demux_001_src6_data),                                               //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src6_startofpacket),                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src6_endofpacket),                                        //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src6_channel),                                            //                .channel
		.rf_sink_ready           (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                      //     (terminated)
		.m0_writeresponserequest (),                                                                           //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                        //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                         // clk_reset.reset
		.in_data           (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                      // (terminated)
		.csr_read          (1'b0),                                                                       // (terminated)
		.csr_write         (1'b0),                                                                       // (terminated)
		.csr_readdata      (),                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                       // (terminated)
		.almost_full_data  (),                                                                           // (terminated)
		.almost_empty_data (),                                                                           // (terminated)
		.in_empty          (1'b0),                                                                       // (terminated)
		.out_empty         (),                                                                           // (terminated)
		.in_error          (1'b0),                                                                       // (terminated)
		.out_error         (),                                                                           // (terminated)
		.in_channel        (1'b0),                                                                       // (terminated)
		.out_channel       ()                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) timer_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                               //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                            //       clk_reset.reset
		.m0_address              (timer_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src7_ready),                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src7_valid),                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_001_src7_data),                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src7_startofpacket),                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src7_endofpacket),                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src7_channel),                                               //                .channel
		.rf_sink_ready           (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                               //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.in_data           (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) performance_counter_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                                        //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                                     //       clk_reset.reset
		.m0_address              (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src8_ready),                                                                          //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src8_valid),                                                                          //                .valid
		.cp_data                 (cmd_xbar_demux_001_src8_data),                                                                           //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src8_startofpacket),                                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src8_endofpacket),                                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src8_channel),                                                                        //                .channel
		.rf_sink_ready           (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                  //     (terminated)
		.m0_writeresponserequest (),                                                                                                       //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                    //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                                        //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                                     // clk_reset.reset
		.in_data           (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                                   // (terminated)
		.csr_readdata      (),                                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                   // (terminated)
		.almost_full_data  (),                                                                                                       // (terminated)
		.almost_empty_data (),                                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                                   // (terminated)
		.out_empty         (),                                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                                   // (terminated)
		.out_error         (),                                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                                   // (terminated)
		.out_channel       ()                                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                              //       clk_reset.reset
		.m0_address              (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src9_ready),                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src9_valid),                                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src9_data),                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src9_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src9_endofpacket),                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src9_channel),                                                                 //                .channel
		.rf_sink_ready           (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                              // clk_reset.reset
		.in_data           (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                           // (terminated)
		.csr_read          (1'b0),                                                                                            // (terminated)
		.csr_write         (1'b0),                                                                                            // (terminated)
		.csr_readdata      (),                                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                            // (terminated)
		.almost_full_data  (),                                                                                                // (terminated)
		.almost_empty_data (),                                                                                                // (terminated)
		.in_empty          (1'b0),                                                                                            // (terminated)
		.out_empty         (),                                                                                                // (terminated)
		.in_error          (1'b0),                                                                                            // (terminated)
		.out_error         (),                                                                                                // (terminated)
		.in_channel        (1'b0),                                                                                            // (terminated)
		.out_channel       ()                                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                              //       clk_reset.reset
		.m0_address              (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src10_ready),                                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src10_valid),                                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src10_data),                                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src10_startofpacket),                                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src10_endofpacket),                                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src10_channel),                                                                //                .channel
		.rf_sink_ready           (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                              // clk_reset.reset
		.in_data           (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                           // (terminated)
		.csr_read          (1'b0),                                                                                            // (terminated)
		.csr_write         (1'b0),                                                                                            // (terminated)
		.csr_readdata      (),                                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                            // (terminated)
		.almost_full_data  (),                                                                                                // (terminated)
		.almost_empty_data (),                                                                                                // (terminated)
		.in_empty          (1'b0),                                                                                            // (terminated)
		.out_empty         (),                                                                                                // (terminated)
		.in_error          (1'b0),                                                                                            // (terminated)
		.out_error         (),                                                                                                // (terminated)
		.in_channel        (1'b0),                                                                                            // (terminated)
		.out_channel       ()                                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) adc_spi_read_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c2_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                      //       clk_reset.reset
		.m0_address              (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_out_ready),                                                                       //              cp.ready
		.cp_valid                (crosser_out_valid),                                                                       //                .valid
		.cp_data                 (crosser_out_data),                                                                        //                .data
		.cp_startofpacket        (crosser_out_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (crosser_out_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (crosser_out_channel),                                                                     //                .channel
		.rf_sink_ready           (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                   //     (terminated)
		.m0_writeresponserequest (),                                                                                        //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                     //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c2_clk),                                                                         //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                      // clk_reset.reset
		.in_data           (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c2_clk),                                                                   //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                // clk_reset.reset
		.in_data           (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_startofpacket  (1'b0),                                                                              // (terminated)
		.in_endofpacket    (1'b0),                                                                              // (terminated)
		.out_startofpacket (),                                                                                  // (terminated)
		.out_endofpacket   (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) pwm0_avalon_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src12_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src12_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_001_src12_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src12_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src12_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src12_channel),                                                       //                .channel
		.rf_sink_ready           (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                  //     (terminated)
		.m0_writeresponserequest (),                                                                                       //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                    //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                        //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) pwm1_avalon_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src13_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src13_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_001_src13_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src13_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src13_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src13_channel),                                                       //                .channel
		.rf_sink_ready           (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                  //     (terminated)
		.m0_writeresponserequest (),                                                                                       //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                    //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                        //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                                    //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                                 //       clk_reset.reset
		.m0_address              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src14_ready),                                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src14_valid),                                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src14_data),                                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src14_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src14_endofpacket),                                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src14_channel),                                                                   //                .channel
		.rf_sink_ready           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                                 // clk_reset.reset
		.in_data           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                              //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src15_ready),                                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src15_valid),                                                               //                .valid
		.cp_data                 (cmd_xbar_demux_001_src15_data),                                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src15_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src15_endofpacket),                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src15_channel),                                                             //                .channel
		.rf_sink_ready           (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                              //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                              //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src16_ready),                                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src16_valid),                                                               //                .valid
		.cp_data                 (cmd_xbar_demux_001_src16_data),                                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src16_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src16_endofpacket),                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src16_channel),                                                             //                .channel
		.rf_sink_ready           (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                              //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) pio_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                               //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                            //       clk_reset.reset
		.m0_address              (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src17_ready),                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src17_valid),                                                //                .valid
		.cp_data                 (cmd_xbar_demux_001_src17_data),                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src17_startofpacket),                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src17_endofpacket),                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src17_channel),                                              //                .channel
		.rf_sink_ready           (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                               //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.in_data           (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) uart_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src18_ready),                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src18_valid),                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_001_src18_data),                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src18_startofpacket),                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src18_endofpacket),                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src18_channel),                                               //                .channel
		.rf_sink_ready           (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                  //       clk_reset.reset
		.m0_address              (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src19_ready),                                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src19_valid),                                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src19_data),                                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src19_startofpacket),                                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src19_endofpacket),                                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src19_channel),                                                                //                .channel
		.rf_sink_ready           (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                  // clk_reset.reset
		.in_data           (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                           // (terminated)
		.csr_read          (1'b0),                                                                                            // (terminated)
		.csr_write         (1'b0),                                                                                            // (terminated)
		.csr_readdata      (),                                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                            // (terminated)
		.almost_full_data  (),                                                                                                // (terminated)
		.almost_empty_data (),                                                                                                // (terminated)
		.in_empty          (1'b0),                                                                                            // (terminated)
		.out_empty         (),                                                                                                // (terminated)
		.in_error          (1'b0),                                                                                            // (terminated)
		.out_error         (),                                                                                                // (terminated)
		.in_channel        (1'b0),                                                                                            // (terminated)
		.out_channel       ()                                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                  //       clk_reset.reset
		.m0_address              (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src20_ready),                                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src20_valid),                                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src20_data),                                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src20_startofpacket),                                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src20_endofpacket),                                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src20_channel),                                                                //                .channel
		.rf_sink_ready           (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                  // clk_reset.reset
		.in_data           (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                           // (terminated)
		.csr_read          (1'b0),                                                                                            // (terminated)
		.csr_write         (1'b0),                                                                                            // (terminated)
		.csr_readdata      (),                                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                            // (terminated)
		.almost_full_data  (),                                                                                                // (terminated)
		.almost_empty_data (),                                                                                                // (terminated)
		.in_empty          (1'b0),                                                                                            // (terminated)
		.out_empty         (),                                                                                                // (terminated)
		.in_error          (1'b0),                                                                                            // (terminated)
		.out_error         (),                                                                                                // (terminated)
		.in_channel        (1'b0),                                                                                            // (terminated)
		.out_channel       ()                                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                  //       clk_reset.reset
		.m0_address              (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src21_ready),                                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src21_valid),                                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src21_data),                                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src21_startofpacket),                                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src21_endofpacket),                                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src21_channel),                                                                //                .channel
		.rf_sink_ready           (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                  // clk_reset.reset
		.in_data           (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                           // (terminated)
		.csr_read          (1'b0),                                                                                            // (terminated)
		.csr_write         (1'b0),                                                                                            // (terminated)
		.csr_readdata      (),                                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                            // (terminated)
		.almost_full_data  (),                                                                                                // (terminated)
		.almost_empty_data (),                                                                                                // (terminated)
		.in_empty          (1'b0),                                                                                            // (terminated)
		.out_empty         (),                                                                                                // (terminated)
		.in_error          (1'b0),                                                                                            // (terminated)
		.out_error         (),                                                                                                // (terminated)
		.in_channel        (1'b0),                                                                                            // (terminated)
		.out_channel       ()                                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                  //       clk_reset.reset
		.m0_address              (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src22_ready),                                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src22_valid),                                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src22_data),                                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src22_startofpacket),                                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src22_endofpacket),                                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src22_channel),                                                                //                .channel
		.rf_sink_ready           (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                  // clk_reset.reset
		.in_data           (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                           // (terminated)
		.csr_read          (1'b0),                                                                                            // (terminated)
		.csr_write         (1'b0),                                                                                            // (terminated)
		.csr_readdata      (),                                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                            // (terminated)
		.almost_full_data  (),                                                                                                // (terminated)
		.almost_empty_data (),                                                                                                // (terminated)
		.in_empty          (1'b0),                                                                                            // (terminated)
		.out_empty         (),                                                                                                // (terminated)
		.in_error          (1'b0),                                                                                            // (terminated)
		.out_error         (),                                                                                                // (terminated)
		.in_channel        (1'b0),                                                                                            // (terminated)
		.out_channel       ()                                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) pwm2_avalon_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src23_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src23_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_001_src23_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src23_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src23_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src23_channel),                                                       //                .channel
		.rf_sink_ready           (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                  //     (terminated)
		.m0_writeresponserequest (),                                                                                       //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                    //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) pwm3_avalon_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src24_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src24_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_001_src24_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src24_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src24_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src24_channel),                                                       //                .channel
		.rf_sink_ready           (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                  //     (terminated)
		.m0_writeresponserequest (),                                                                                       //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                    //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) pio_1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pio_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pio_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pio_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pio_1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pio_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src25_ready),                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src25_valid),                                                //                .valid
		.cp_data                 (cmd_xbar_demux_001_src25_data),                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src25_startofpacket),                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src25_endofpacket),                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src25_channel),                                              //                .channel
		.rf_sink_ready           (pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.in_data           (pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	NIOS_Sys_addr_router addr_router (
		.sink_ready         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                       //       src.ready
		.src_valid          (addr_router_src_valid),                                                                       //          .valid
		.src_data           (addr_router_src_data),                                                                        //          .data
		.src_channel        (addr_router_src_channel),                                                                     //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                               //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                                  //          .endofpacket
	);

	NIOS_Sys_addr_router_001 addr_router_001 (
		.sink_ready         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                            //          .valid
		.src_data           (addr_router_001_src_data),                                                             //          .data
		.src_channel        (addr_router_001_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                       //          .endofpacket
	);

	NIOS_Sys_id_router id_router (
		.sink_ready         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                       //       src.ready
		.src_valid          (id_router_src_valid),                                                                       //          .valid
		.src_data           (id_router_src_data),                                                                        //          .data
		.src_channel        (id_router_src_channel),                                                                     //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                               //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                                  //          .endofpacket
	);

	NIOS_Sys_id_router_001 id_router_001 (
		.sink_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                     //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                  // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                             //       src.ready
		.src_valid          (id_router_001_src_valid),                                             //          .valid
		.src_data           (id_router_001_src_data),                                              //          .data
		.src_channel        (id_router_001_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                        //          .endofpacket
	);

	NIOS_Sys_id_router id_router_002 (
		.sink_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                        //       src.ready
		.src_valid          (id_router_002_src_valid),                                                        //          .valid
		.src_data           (id_router_002_src_data),                                                         //          .data
		.src_channel        (id_router_002_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                   //          .endofpacket
	);

	NIOS_Sys_id_router id_router_003 (
		.sink_ready         (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                       // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                                              //       src.ready
		.src_valid          (id_router_003_src_valid),                                                                              //          .valid
		.src_data           (id_router_003_src_data),                                                                               //          .data
		.src_channel        (id_router_003_src_channel),                                                                            //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                                      //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                                         //          .endofpacket
	);

	NIOS_Sys_id_router_004 id_router_004 (
		.sink_ready         (led_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (led_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (led_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                           //       src.ready
		.src_valid          (id_router_004_src_valid),                                           //          .valid
		.src_data           (id_router_004_src_data),                                            //          .data
		.src_channel        (id_router_004_src_channel),                                         //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                   //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                      //          .endofpacket
	);

	NIOS_Sys_id_router_004 id_router_005 (
		.sink_ready         (key_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (key_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (key_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (key_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (key_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                           //       src.ready
		.src_valid          (id_router_005_src_valid),                                           //          .valid
		.src_data           (id_router_005_src_data),                                            //          .data
		.src_channel        (id_router_005_src_channel),                                         //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                   //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                      //          .endofpacket
	);

	NIOS_Sys_id_router_004 id_router_006 (
		.sink_ready         (sw_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sw_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sw_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                               // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                          //       src.ready
		.src_valid          (id_router_006_src_valid),                                          //          .valid
		.src_data           (id_router_006_src_data),                                           //          .data
		.src_channel        (id_router_006_src_channel),                                        //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                  //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                     //          .endofpacket
	);

	NIOS_Sys_id_router_004 id_router_007 (
		.sink_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                     //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                  // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                             //       src.ready
		.src_valid          (id_router_007_src_valid),                                             //          .valid
		.src_data           (id_router_007_src_data),                                              //          .data
		.src_channel        (id_router_007_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                        //          .endofpacket
	);

	NIOS_Sys_id_router_004 id_router_008 (
		.sink_ready         (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                              //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                                      //       src.ready
		.src_valid          (id_router_008_src_valid),                                                                      //          .valid
		.src_data           (id_router_008_src_data),                                                                       //          .data
		.src_channel        (id_router_008_src_channel),                                                                    //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                                              //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                                                 //          .endofpacket
	);

	NIOS_Sys_id_router_004 id_router_009 (
		.sink_ready         (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ultrasound0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                                               //       src.ready
		.src_valid          (id_router_009_src_valid),                                                               //          .valid
		.src_data           (id_router_009_src_data),                                                                //          .data
		.src_channel        (id_router_009_src_channel),                                                             //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                                       //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                                          //          .endofpacket
	);

	NIOS_Sys_id_router_004 id_router_010 (
		.sink_ready         (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ultrasound1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                                               //       src.ready
		.src_valid          (id_router_010_src_valid),                                                               //          .valid
		.src_data           (id_router_010_src_data),                                                                //          .data
		.src_channel        (id_router_010_src_channel),                                                             //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                                       //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                                          //          .endofpacket
	);

	NIOS_Sys_id_router_004 id_router_011 (
		.sink_ready         (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (adc_spi_read_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c2_clk),                                                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                            // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                                       //       src.ready
		.src_valid          (id_router_011_src_valid),                                                       //          .valid
		.src_data           (id_router_011_src_data),                                                        //          .data
		.src_channel        (id_router_011_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                                  //          .endofpacket
	);

	NIOS_Sys_id_router_004 id_router_012 (
		.sink_ready         (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pwm0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                              //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                                      //       src.ready
		.src_valid          (id_router_012_src_valid),                                                      //          .valid
		.src_data           (id_router_012_src_data),                                                       //          .data
		.src_channel        (id_router_012_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                                 //          .endofpacket
	);

	NIOS_Sys_id_router_004 id_router_013 (
		.sink_ready         (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pwm1_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                              //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                                      //       src.ready
		.src_valid          (id_router_013_src_valid),                                                      //          .valid
		.src_data           (id_router_013_src_data),                                                       //          .data
		.src_channel        (id_router_013_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                                 //          .endofpacket
	);

	NIOS_Sys_id_router_004 id_router_014 (
		.sink_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                          //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (id_router_014_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_014_src_valid),                                                                  //          .valid
		.src_data           (id_router_014_src_data),                                                                   //          .data
		.src_channel        (id_router_014_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_014_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_014_src_endofpacket)                                                             //          .endofpacket
	);

	NIOS_Sys_id_router_004 id_router_015 (
		.sink_ready         (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (encoder0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                    //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_015_src_ready),                                                            //       src.ready
		.src_valid          (id_router_015_src_valid),                                                            //          .valid
		.src_data           (id_router_015_src_data),                                                             //          .data
		.src_channel        (id_router_015_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_015_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_015_src_endofpacket)                                                       //          .endofpacket
	);

	NIOS_Sys_id_router_004 id_router_016 (
		.sink_ready         (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (encoder1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                    //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_016_src_ready),                                                            //       src.ready
		.src_valid          (id_router_016_src_valid),                                                            //          .valid
		.src_data           (id_router_016_src_data),                                                             //          .data
		.src_channel        (id_router_016_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_016_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_016_src_endofpacket)                                                       //          .endofpacket
	);

	NIOS_Sys_id_router_004 id_router_017 (
		.sink_ready         (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                     //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                  // clk_reset.reset
		.src_ready          (id_router_017_src_ready),                                             //       src.ready
		.src_valid          (id_router_017_src_valid),                                             //          .valid
		.src_data           (id_router_017_src_data),                                              //          .data
		.src_channel        (id_router_017_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_017_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_017_src_endofpacket)                                        //          .endofpacket
	);

	NIOS_Sys_id_router_004 id_router_018 (
		.sink_ready         (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_018_src_ready),                                              //       src.ready
		.src_valid          (id_router_018_src_valid),                                              //          .valid
		.src_data           (id_router_018_src_data),                                               //          .data
		.src_channel        (id_router_018_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_018_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_018_src_endofpacket)                                         //          .endofpacket
	);

	NIOS_Sys_id_router_004 id_router_019 (
		.sink_ready         (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ultrasound2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.src_ready          (id_router_019_src_ready),                                                               //       src.ready
		.src_valid          (id_router_019_src_valid),                                                               //          .valid
		.src_data           (id_router_019_src_data),                                                                //          .data
		.src_channel        (id_router_019_src_channel),                                                             //          .channel
		.src_startofpacket  (id_router_019_src_startofpacket),                                                       //          .startofpacket
		.src_endofpacket    (id_router_019_src_endofpacket)                                                          //          .endofpacket
	);

	NIOS_Sys_id_router_004 id_router_020 (
		.sink_ready         (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ultrasound3_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.src_ready          (id_router_020_src_ready),                                                               //       src.ready
		.src_valid          (id_router_020_src_valid),                                                               //          .valid
		.src_data           (id_router_020_src_data),                                                                //          .data
		.src_channel        (id_router_020_src_channel),                                                             //          .channel
		.src_startofpacket  (id_router_020_src_startofpacket),                                                       //          .startofpacket
		.src_endofpacket    (id_router_020_src_endofpacket)                                                          //          .endofpacket
	);

	NIOS_Sys_id_router_004 id_router_021 (
		.sink_ready         (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ultrasound4_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.src_ready          (id_router_021_src_ready),                                                               //       src.ready
		.src_valid          (id_router_021_src_valid),                                                               //          .valid
		.src_data           (id_router_021_src_data),                                                                //          .data
		.src_channel        (id_router_021_src_channel),                                                             //          .channel
		.src_startofpacket  (id_router_021_src_startofpacket),                                                       //          .startofpacket
		.src_endofpacket    (id_router_021_src_endofpacket)                                                          //          .endofpacket
	);

	NIOS_Sys_id_router_004 id_router_022 (
		.sink_ready         (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ultrasound5_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.src_ready          (id_router_022_src_ready),                                                               //       src.ready
		.src_valid          (id_router_022_src_valid),                                                               //          .valid
		.src_data           (id_router_022_src_data),                                                                //          .data
		.src_channel        (id_router_022_src_channel),                                                             //          .channel
		.src_startofpacket  (id_router_022_src_startofpacket),                                                       //          .startofpacket
		.src_endofpacket    (id_router_022_src_endofpacket)                                                          //          .endofpacket
	);

	NIOS_Sys_id_router_004 id_router_023 (
		.sink_ready         (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pwm2_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_023_src_ready),                                                      //       src.ready
		.src_valid          (id_router_023_src_valid),                                                      //          .valid
		.src_data           (id_router_023_src_data),                                                       //          .data
		.src_channel        (id_router_023_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_023_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_023_src_endofpacket)                                                 //          .endofpacket
	);

	NIOS_Sys_id_router_004 id_router_024 (
		.sink_ready         (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pwm3_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_024_src_ready),                                                      //       src.ready
		.src_valid          (id_router_024_src_valid),                                                      //          .valid
		.src_data           (id_router_024_src_data),                                                       //          .data
		.src_channel        (id_router_024_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_024_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_024_src_endofpacket)                                                 //          .endofpacket
	);

	NIOS_Sys_id_router_004 id_router_025 (
		.sink_ready         (pio_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pio_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pio_1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pio_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pio_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_025_src_ready),                                             //       src.ready
		.src_valid          (id_router_025_src_valid),                                             //          .valid
		.src_data           (id_router_025_src_data),                                              //          .data
		.src_channel        (id_router_025_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_025_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_025_src_endofpacket)                                        //          .endofpacket
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (43),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (63),
		.PKT_BYTE_CNT_H            (52),
		.PKT_BYTE_CNT_L            (50),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.PKT_BURST_TYPE_H          (60),
		.PKT_BURST_TYPE_L          (59),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (53),
		.PKT_TRANS_COMPRESSED_READ (44),
		.PKT_TRANS_WRITE           (46),
		.PKT_TRANS_READ            (47),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (85),
		.ST_CHANNEL_W              (26),
		.OUT_BYTE_CNT_H            (51),
		.OUT_BURSTWRAP_H           (55),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter (
		.clk                   (altpll_0_c0_clk),                     //       cr0.clk
		.reset                 (rst_controller_001_reset_out_reset),  // cr0_reset.reset
		.sink0_valid           (width_adapter_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_src_data),              //          .data
		.sink0_channel         (width_adapter_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_src_ready),             //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (altpll_0_c0_clk),                //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req  (),                               // (terminated)
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (1)
	) rst_controller_001 (
		.reset_in0  (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1  (~reset_reset_n),                             // reset_in1.reset
		.clk        (altpll_0_c0_clk),                            //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset),         // reset_out.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),     //          .reset_req
		.reset_in2  (1'b0),                                       // (terminated)
		.reset_in3  (1'b0),                                       // (terminated)
		.reset_in4  (1'b0),                                       // (terminated)
		.reset_in5  (1'b0),                                       // (terminated)
		.reset_in6  (1'b0),                                       // (terminated)
		.reset_in7  (1'b0),                                       // (terminated)
		.reset_in8  (1'b0),                                       // (terminated)
		.reset_in9  (1'b0),                                       // (terminated)
		.reset_in10 (1'b0),                                       // (terminated)
		.reset_in11 (1'b0),                                       // (terminated)
		.reset_in12 (1'b0),                                       // (terminated)
		.reset_in13 (1'b0),                                       // (terminated)
		.reset_in14 (1'b0),                                       // (terminated)
		.reset_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_002 (
		.reset_in0  (~reset_reset_n),                             // reset_in0.reset
		.reset_in1  (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_clk),                                    //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset),         // reset_out.reset
		.reset_req  (),                                           // (terminated)
		.reset_in2  (1'b0),                                       // (terminated)
		.reset_in3  (1'b0),                                       // (terminated)
		.reset_in4  (1'b0),                                       // (terminated)
		.reset_in5  (1'b0),                                       // (terminated)
		.reset_in6  (1'b0),                                       // (terminated)
		.reset_in7  (1'b0),                                       // (terminated)
		.reset_in8  (1'b0),                                       // (terminated)
		.reset_in9  (1'b0),                                       // (terminated)
		.reset_in10 (1'b0),                                       // (terminated)
		.reset_in11 (1'b0),                                       // (terminated)
		.reset_in12 (1'b0),                                       // (terminated)
		.reset_in13 (1'b0),                                       // (terminated)
		.reset_in14 (1'b0),                                       // (terminated)
		.reset_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_003 (
		.reset_in0  (~reset_reset_n),                             // reset_in0.reset
		.reset_in1  (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (altpll_0_c2_clk),                            //       clk.clk
		.reset_out  (rst_controller_003_reset_out_reset),         // reset_out.reset
		.reset_req  (),                                           // (terminated)
		.reset_in2  (1'b0),                                       // (terminated)
		.reset_in3  (1'b0),                                       // (terminated)
		.reset_in4  (1'b0),                                       // (terminated)
		.reset_in5  (1'b0),                                       // (terminated)
		.reset_in6  (1'b0),                                       // (terminated)
		.reset_in7  (1'b0),                                       // (terminated)
		.reset_in8  (1'b0),                                       // (terminated)
		.reset_in9  (1'b0),                                       // (terminated)
		.reset_in10 (1'b0),                                       // (terminated)
		.reset_in11 (1'b0),                                       // (terminated)
		.reset_in12 (1'b0),                                       // (terminated)
		.reset_in13 (1'b0),                                       // (terminated)
		.reset_in14 (1'b0),                                       // (terminated)
		.reset_in15 (1'b0)                                        // (terminated)
	);

	NIOS_Sys_cmd_xbar_demux cmd_xbar_demux (
		.clk                (altpll_0_c0_clk),                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_src_ready),             //      sink.ready
		.sink_channel       (addr_router_src_channel),           //          .channel
		.sink_data          (addr_router_src_data),              //          .data
		.sink_startofpacket (addr_router_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),   //          .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),         //      src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),         //          .valid
		.src2_data          (cmd_xbar_demux_src2_data),          //          .data
		.src2_channel       (cmd_xbar_demux_src2_channel),       //          .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket),   //          .endofpacket
		.src3_ready         (cmd_xbar_demux_src3_ready),         //      src3.ready
		.src3_valid         (cmd_xbar_demux_src3_valid),         //          .valid
		.src3_data          (cmd_xbar_demux_src3_data),          //          .data
		.src3_channel       (cmd_xbar_demux_src3_channel),       //          .channel
		.src3_startofpacket (cmd_xbar_demux_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_src3_endofpacket)    //          .endofpacket
	);

	NIOS_Sys_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                 (altpll_0_c0_clk),                        //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.sink_ready          (addr_router_001_src_ready),              //      sink.ready
		.sink_channel        (addr_router_001_src_channel),            //          .channel
		.sink_data           (addr_router_001_src_data),               //          .data
		.sink_startofpacket  (addr_router_001_src_startofpacket),      //          .startofpacket
		.sink_endofpacket    (addr_router_001_src_endofpacket),        //          .endofpacket
		.sink_valid          (addr_router_001_src_valid),              //          .valid
		.src0_ready          (cmd_xbar_demux_001_src0_ready),          //      src0.ready
		.src0_valid          (cmd_xbar_demux_001_src0_valid),          //          .valid
		.src0_data           (cmd_xbar_demux_001_src0_data),           //          .data
		.src0_channel        (cmd_xbar_demux_001_src0_channel),        //          .channel
		.src0_startofpacket  (cmd_xbar_demux_001_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_001_src0_endofpacket),    //          .endofpacket
		.src1_ready          (cmd_xbar_demux_001_src1_ready),          //      src1.ready
		.src1_valid          (cmd_xbar_demux_001_src1_valid),          //          .valid
		.src1_data           (cmd_xbar_demux_001_src1_data),           //          .data
		.src1_channel        (cmd_xbar_demux_001_src1_channel),        //          .channel
		.src1_startofpacket  (cmd_xbar_demux_001_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_001_src1_endofpacket),    //          .endofpacket
		.src2_ready          (cmd_xbar_demux_001_src2_ready),          //      src2.ready
		.src2_valid          (cmd_xbar_demux_001_src2_valid),          //          .valid
		.src2_data           (cmd_xbar_demux_001_src2_data),           //          .data
		.src2_channel        (cmd_xbar_demux_001_src2_channel),        //          .channel
		.src2_startofpacket  (cmd_xbar_demux_001_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_001_src2_endofpacket),    //          .endofpacket
		.src3_ready          (cmd_xbar_demux_001_src3_ready),          //      src3.ready
		.src3_valid          (cmd_xbar_demux_001_src3_valid),          //          .valid
		.src3_data           (cmd_xbar_demux_001_src3_data),           //          .data
		.src3_channel        (cmd_xbar_demux_001_src3_channel),        //          .channel
		.src3_startofpacket  (cmd_xbar_demux_001_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_001_src3_endofpacket),    //          .endofpacket
		.src4_ready          (cmd_xbar_demux_001_src4_ready),          //      src4.ready
		.src4_valid          (cmd_xbar_demux_001_src4_valid),          //          .valid
		.src4_data           (cmd_xbar_demux_001_src4_data),           //          .data
		.src4_channel        (cmd_xbar_demux_001_src4_channel),        //          .channel
		.src4_startofpacket  (cmd_xbar_demux_001_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_001_src4_endofpacket),    //          .endofpacket
		.src5_ready          (cmd_xbar_demux_001_src5_ready),          //      src5.ready
		.src5_valid          (cmd_xbar_demux_001_src5_valid),          //          .valid
		.src5_data           (cmd_xbar_demux_001_src5_data),           //          .data
		.src5_channel        (cmd_xbar_demux_001_src5_channel),        //          .channel
		.src5_startofpacket  (cmd_xbar_demux_001_src5_startofpacket),  //          .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_001_src5_endofpacket),    //          .endofpacket
		.src6_ready          (cmd_xbar_demux_001_src6_ready),          //      src6.ready
		.src6_valid          (cmd_xbar_demux_001_src6_valid),          //          .valid
		.src6_data           (cmd_xbar_demux_001_src6_data),           //          .data
		.src6_channel        (cmd_xbar_demux_001_src6_channel),        //          .channel
		.src6_startofpacket  (cmd_xbar_demux_001_src6_startofpacket),  //          .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_001_src6_endofpacket),    //          .endofpacket
		.src7_ready          (cmd_xbar_demux_001_src7_ready),          //      src7.ready
		.src7_valid          (cmd_xbar_demux_001_src7_valid),          //          .valid
		.src7_data           (cmd_xbar_demux_001_src7_data),           //          .data
		.src7_channel        (cmd_xbar_demux_001_src7_channel),        //          .channel
		.src7_startofpacket  (cmd_xbar_demux_001_src7_startofpacket),  //          .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_001_src7_endofpacket),    //          .endofpacket
		.src8_ready          (cmd_xbar_demux_001_src8_ready),          //      src8.ready
		.src8_valid          (cmd_xbar_demux_001_src8_valid),          //          .valid
		.src8_data           (cmd_xbar_demux_001_src8_data),           //          .data
		.src8_channel        (cmd_xbar_demux_001_src8_channel),        //          .channel
		.src8_startofpacket  (cmd_xbar_demux_001_src8_startofpacket),  //          .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_001_src8_endofpacket),    //          .endofpacket
		.src9_ready          (cmd_xbar_demux_001_src9_ready),          //      src9.ready
		.src9_valid          (cmd_xbar_demux_001_src9_valid),          //          .valid
		.src9_data           (cmd_xbar_demux_001_src9_data),           //          .data
		.src9_channel        (cmd_xbar_demux_001_src9_channel),        //          .channel
		.src9_startofpacket  (cmd_xbar_demux_001_src9_startofpacket),  //          .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_001_src9_endofpacket),    //          .endofpacket
		.src10_ready         (cmd_xbar_demux_001_src10_ready),         //     src10.ready
		.src10_valid         (cmd_xbar_demux_001_src10_valid),         //          .valid
		.src10_data          (cmd_xbar_demux_001_src10_data),          //          .data
		.src10_channel       (cmd_xbar_demux_001_src10_channel),       //          .channel
		.src10_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //          .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_001_src10_endofpacket),   //          .endofpacket
		.src11_ready         (cmd_xbar_demux_001_src11_ready),         //     src11.ready
		.src11_valid         (cmd_xbar_demux_001_src11_valid),         //          .valid
		.src11_data          (cmd_xbar_demux_001_src11_data),          //          .data
		.src11_channel       (cmd_xbar_demux_001_src11_channel),       //          .channel
		.src11_startofpacket (cmd_xbar_demux_001_src11_startofpacket), //          .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_001_src11_endofpacket),   //          .endofpacket
		.src12_ready         (cmd_xbar_demux_001_src12_ready),         //     src12.ready
		.src12_valid         (cmd_xbar_demux_001_src12_valid),         //          .valid
		.src12_data          (cmd_xbar_demux_001_src12_data),          //          .data
		.src12_channel       (cmd_xbar_demux_001_src12_channel),       //          .channel
		.src12_startofpacket (cmd_xbar_demux_001_src12_startofpacket), //          .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_001_src12_endofpacket),   //          .endofpacket
		.src13_ready         (cmd_xbar_demux_001_src13_ready),         //     src13.ready
		.src13_valid         (cmd_xbar_demux_001_src13_valid),         //          .valid
		.src13_data          (cmd_xbar_demux_001_src13_data),          //          .data
		.src13_channel       (cmd_xbar_demux_001_src13_channel),       //          .channel
		.src13_startofpacket (cmd_xbar_demux_001_src13_startofpacket), //          .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_001_src13_endofpacket),   //          .endofpacket
		.src14_ready         (cmd_xbar_demux_001_src14_ready),         //     src14.ready
		.src14_valid         (cmd_xbar_demux_001_src14_valid),         //          .valid
		.src14_data          (cmd_xbar_demux_001_src14_data),          //          .data
		.src14_channel       (cmd_xbar_demux_001_src14_channel),       //          .channel
		.src14_startofpacket (cmd_xbar_demux_001_src14_startofpacket), //          .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_001_src14_endofpacket),   //          .endofpacket
		.src15_ready         (cmd_xbar_demux_001_src15_ready),         //     src15.ready
		.src15_valid         (cmd_xbar_demux_001_src15_valid),         //          .valid
		.src15_data          (cmd_xbar_demux_001_src15_data),          //          .data
		.src15_channel       (cmd_xbar_demux_001_src15_channel),       //          .channel
		.src15_startofpacket (cmd_xbar_demux_001_src15_startofpacket), //          .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_001_src15_endofpacket),   //          .endofpacket
		.src16_ready         (cmd_xbar_demux_001_src16_ready),         //     src16.ready
		.src16_valid         (cmd_xbar_demux_001_src16_valid),         //          .valid
		.src16_data          (cmd_xbar_demux_001_src16_data),          //          .data
		.src16_channel       (cmd_xbar_demux_001_src16_channel),       //          .channel
		.src16_startofpacket (cmd_xbar_demux_001_src16_startofpacket), //          .startofpacket
		.src16_endofpacket   (cmd_xbar_demux_001_src16_endofpacket),   //          .endofpacket
		.src17_ready         (cmd_xbar_demux_001_src17_ready),         //     src17.ready
		.src17_valid         (cmd_xbar_demux_001_src17_valid),         //          .valid
		.src17_data          (cmd_xbar_demux_001_src17_data),          //          .data
		.src17_channel       (cmd_xbar_demux_001_src17_channel),       //          .channel
		.src17_startofpacket (cmd_xbar_demux_001_src17_startofpacket), //          .startofpacket
		.src17_endofpacket   (cmd_xbar_demux_001_src17_endofpacket),   //          .endofpacket
		.src18_ready         (cmd_xbar_demux_001_src18_ready),         //     src18.ready
		.src18_valid         (cmd_xbar_demux_001_src18_valid),         //          .valid
		.src18_data          (cmd_xbar_demux_001_src18_data),          //          .data
		.src18_channel       (cmd_xbar_demux_001_src18_channel),       //          .channel
		.src18_startofpacket (cmd_xbar_demux_001_src18_startofpacket), //          .startofpacket
		.src18_endofpacket   (cmd_xbar_demux_001_src18_endofpacket),   //          .endofpacket
		.src19_ready         (cmd_xbar_demux_001_src19_ready),         //     src19.ready
		.src19_valid         (cmd_xbar_demux_001_src19_valid),         //          .valid
		.src19_data          (cmd_xbar_demux_001_src19_data),          //          .data
		.src19_channel       (cmd_xbar_demux_001_src19_channel),       //          .channel
		.src19_startofpacket (cmd_xbar_demux_001_src19_startofpacket), //          .startofpacket
		.src19_endofpacket   (cmd_xbar_demux_001_src19_endofpacket),   //          .endofpacket
		.src20_ready         (cmd_xbar_demux_001_src20_ready),         //     src20.ready
		.src20_valid         (cmd_xbar_demux_001_src20_valid),         //          .valid
		.src20_data          (cmd_xbar_demux_001_src20_data),          //          .data
		.src20_channel       (cmd_xbar_demux_001_src20_channel),       //          .channel
		.src20_startofpacket (cmd_xbar_demux_001_src20_startofpacket), //          .startofpacket
		.src20_endofpacket   (cmd_xbar_demux_001_src20_endofpacket),   //          .endofpacket
		.src21_ready         (cmd_xbar_demux_001_src21_ready),         //     src21.ready
		.src21_valid         (cmd_xbar_demux_001_src21_valid),         //          .valid
		.src21_data          (cmd_xbar_demux_001_src21_data),          //          .data
		.src21_channel       (cmd_xbar_demux_001_src21_channel),       //          .channel
		.src21_startofpacket (cmd_xbar_demux_001_src21_startofpacket), //          .startofpacket
		.src21_endofpacket   (cmd_xbar_demux_001_src21_endofpacket),   //          .endofpacket
		.src22_ready         (cmd_xbar_demux_001_src22_ready),         //     src22.ready
		.src22_valid         (cmd_xbar_demux_001_src22_valid),         //          .valid
		.src22_data          (cmd_xbar_demux_001_src22_data),          //          .data
		.src22_channel       (cmd_xbar_demux_001_src22_channel),       //          .channel
		.src22_startofpacket (cmd_xbar_demux_001_src22_startofpacket), //          .startofpacket
		.src22_endofpacket   (cmd_xbar_demux_001_src22_endofpacket),   //          .endofpacket
		.src23_ready         (cmd_xbar_demux_001_src23_ready),         //     src23.ready
		.src23_valid         (cmd_xbar_demux_001_src23_valid),         //          .valid
		.src23_data          (cmd_xbar_demux_001_src23_data),          //          .data
		.src23_channel       (cmd_xbar_demux_001_src23_channel),       //          .channel
		.src23_startofpacket (cmd_xbar_demux_001_src23_startofpacket), //          .startofpacket
		.src23_endofpacket   (cmd_xbar_demux_001_src23_endofpacket),   //          .endofpacket
		.src24_ready         (cmd_xbar_demux_001_src24_ready),         //     src24.ready
		.src24_valid         (cmd_xbar_demux_001_src24_valid),         //          .valid
		.src24_data          (cmd_xbar_demux_001_src24_data),          //          .data
		.src24_channel       (cmd_xbar_demux_001_src24_channel),       //          .channel
		.src24_startofpacket (cmd_xbar_demux_001_src24_startofpacket), //          .startofpacket
		.src24_endofpacket   (cmd_xbar_demux_001_src24_endofpacket),   //          .endofpacket
		.src25_ready         (cmd_xbar_demux_001_src25_ready),         //     src25.ready
		.src25_valid         (cmd_xbar_demux_001_src25_valid),         //          .valid
		.src25_data          (cmd_xbar_demux_001_src25_data),          //          .data
		.src25_channel       (cmd_xbar_demux_001_src25_channel),       //          .channel
		.src25_startofpacket (cmd_xbar_demux_001_src25_startofpacket), //          .startofpacket
		.src25_endofpacket   (cmd_xbar_demux_001_src25_endofpacket)    //          .endofpacket
	);

	NIOS_Sys_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (altpll_0_c0_clk),                       //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	NIOS_Sys_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (altpll_0_c0_clk),                       //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	NIOS_Sys_cmd_xbar_mux cmd_xbar_mux_002 (
		.clk                 (altpll_0_c0_clk),                       //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src2_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src2_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src2_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src2_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src2_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src2_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)    //          .endofpacket
	);

	NIOS_Sys_cmd_xbar_mux cmd_xbar_mux_003 (
		.clk                 (altpll_0_c0_clk),                       //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_003_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_003_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src3_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src3_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src3_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src3_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src3_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src3_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src3_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src3_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src3_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src3_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src3_endofpacket)    //          .endofpacket
	);

	NIOS_Sys_rsp_xbar_demux rsp_xbar_demux (
		.clk                (altpll_0_c0_clk),                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	NIOS_Sys_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (width_adapter_001_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_001_src_channel),         //          .channel
		.sink_data          (width_adapter_001_src_data),            //          .data
		.sink_startofpacket (width_adapter_001_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_001_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_001_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	NIOS_Sys_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	NIOS_Sys_rsp_xbar_demux rsp_xbar_demux_003 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_003_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_003_src1_endofpacket)    //          .endofpacket
	);

	NIOS_Sys_rsp_xbar_demux_004 rsp_xbar_demux_004 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	NIOS_Sys_rsp_xbar_demux_004 rsp_xbar_demux_005 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	NIOS_Sys_rsp_xbar_demux_004 rsp_xbar_demux_006 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	NIOS_Sys_rsp_xbar_demux_004 rsp_xbar_demux_007 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	NIOS_Sys_rsp_xbar_demux_004 rsp_xbar_demux_008 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	NIOS_Sys_rsp_xbar_demux_004 rsp_xbar_demux_009 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	NIOS_Sys_rsp_xbar_demux_004 rsp_xbar_demux_010 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	NIOS_Sys_rsp_xbar_demux_004 rsp_xbar_demux_011 (
		.clk                (altpll_0_c2_clk),                       //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	NIOS_Sys_rsp_xbar_demux_004 rsp_xbar_demux_012 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	NIOS_Sys_rsp_xbar_demux_004 rsp_xbar_demux_013 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket)    //          .endofpacket
	);

	NIOS_Sys_rsp_xbar_demux_004 rsp_xbar_demux_014 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_014_src_ready),               //      sink.ready
		.sink_channel       (id_router_014_src_channel),             //          .channel
		.sink_data          (id_router_014_src_data),                //          .data
		.sink_startofpacket (id_router_014_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_014_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_014_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket)    //          .endofpacket
	);

	NIOS_Sys_rsp_xbar_demux_004 rsp_xbar_demux_015 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_015_src_ready),               //      sink.ready
		.sink_channel       (id_router_015_src_channel),             //          .channel
		.sink_data          (id_router_015_src_data),                //          .data
		.sink_startofpacket (id_router_015_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_015_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_015_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_015_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_015_src0_endofpacket)    //          .endofpacket
	);

	NIOS_Sys_rsp_xbar_demux_004 rsp_xbar_demux_016 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_016_src_ready),               //      sink.ready
		.sink_channel       (id_router_016_src_channel),             //          .channel
		.sink_data          (id_router_016_src_data),                //          .data
		.sink_startofpacket (id_router_016_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_016_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_016_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_016_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_016_src0_endofpacket)    //          .endofpacket
	);

	NIOS_Sys_rsp_xbar_demux_004 rsp_xbar_demux_017 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_017_src_ready),               //      sink.ready
		.sink_channel       (id_router_017_src_channel),             //          .channel
		.sink_data          (id_router_017_src_data),                //          .data
		.sink_startofpacket (id_router_017_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_017_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_017_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_017_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_017_src0_endofpacket)    //          .endofpacket
	);

	NIOS_Sys_rsp_xbar_demux_004 rsp_xbar_demux_018 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_018_src_ready),               //      sink.ready
		.sink_channel       (id_router_018_src_channel),             //          .channel
		.sink_data          (id_router_018_src_data),                //          .data
		.sink_startofpacket (id_router_018_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_018_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_018_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_018_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_018_src0_endofpacket)    //          .endofpacket
	);

	NIOS_Sys_rsp_xbar_demux_004 rsp_xbar_demux_019 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_019_src_ready),               //      sink.ready
		.sink_channel       (id_router_019_src_channel),             //          .channel
		.sink_data          (id_router_019_src_data),                //          .data
		.sink_startofpacket (id_router_019_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_019_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_019_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_019_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_019_src0_endofpacket)    //          .endofpacket
	);

	NIOS_Sys_rsp_xbar_demux_004 rsp_xbar_demux_020 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_020_src_ready),               //      sink.ready
		.sink_channel       (id_router_020_src_channel),             //          .channel
		.sink_data          (id_router_020_src_data),                //          .data
		.sink_startofpacket (id_router_020_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_020_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_020_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_020_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_020_src0_endofpacket)    //          .endofpacket
	);

	NIOS_Sys_rsp_xbar_demux_004 rsp_xbar_demux_021 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_021_src_ready),               //      sink.ready
		.sink_channel       (id_router_021_src_channel),             //          .channel
		.sink_data          (id_router_021_src_data),                //          .data
		.sink_startofpacket (id_router_021_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_021_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_021_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_021_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_021_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_021_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_021_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_021_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_021_src0_endofpacket)    //          .endofpacket
	);

	NIOS_Sys_rsp_xbar_demux_004 rsp_xbar_demux_022 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_022_src_ready),               //      sink.ready
		.sink_channel       (id_router_022_src_channel),             //          .channel
		.sink_data          (id_router_022_src_data),                //          .data
		.sink_startofpacket (id_router_022_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_022_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_022_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_022_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_022_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_022_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_022_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_022_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_022_src0_endofpacket)    //          .endofpacket
	);

	NIOS_Sys_rsp_xbar_demux_004 rsp_xbar_demux_023 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_023_src_ready),               //      sink.ready
		.sink_channel       (id_router_023_src_channel),             //          .channel
		.sink_data          (id_router_023_src_data),                //          .data
		.sink_startofpacket (id_router_023_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_023_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_023_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_023_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_023_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_023_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_023_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_023_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_023_src0_endofpacket)    //          .endofpacket
	);

	NIOS_Sys_rsp_xbar_demux_004 rsp_xbar_demux_024 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_024_src_ready),               //      sink.ready
		.sink_channel       (id_router_024_src_channel),             //          .channel
		.sink_data          (id_router_024_src_data),                //          .data
		.sink_startofpacket (id_router_024_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_024_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_024_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_024_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_024_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_024_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_024_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_024_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_024_src0_endofpacket)    //          .endofpacket
	);

	NIOS_Sys_rsp_xbar_demux_004 rsp_xbar_demux_025 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_025_src_ready),               //      sink.ready
		.sink_channel       (id_router_025_src_channel),             //          .channel
		.sink_data          (id_router_025_src_data),                //          .data
		.sink_startofpacket (id_router_025_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_025_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_025_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_025_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_025_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_025_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_025_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_025_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_025_src0_endofpacket)    //          .endofpacket
	);

	NIOS_Sys_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (altpll_0_c0_clk),                       //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	NIOS_Sys_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                  (altpll_0_c0_clk),                       //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_002_src1_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_002_src1_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_002_src1_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_002_src1_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_003_src1_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_003_src1_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_003_src1_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_003_src1_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_010_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (crosser_001_out_ready),                 //    sink11.ready
		.sink11_valid         (crosser_001_out_valid),                 //          .valid
		.sink11_channel       (crosser_001_out_channel),               //          .channel
		.sink11_data          (crosser_001_out_data),                  //          .data
		.sink11_startofpacket (crosser_001_out_startofpacket),         //          .startofpacket
		.sink11_endofpacket   (crosser_001_out_endofpacket),           //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_012_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_013_src0_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.sink14_ready         (rsp_xbar_demux_014_src0_ready),         //    sink14.ready
		.sink14_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.sink14_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.sink14_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.sink14_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.sink14_endofpacket   (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.sink15_ready         (rsp_xbar_demux_015_src0_ready),         //    sink15.ready
		.sink15_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.sink15_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.sink15_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.sink15_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.sink15_endofpacket   (rsp_xbar_demux_015_src0_endofpacket),   //          .endofpacket
		.sink16_ready         (rsp_xbar_demux_016_src0_ready),         //    sink16.ready
		.sink16_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.sink16_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.sink16_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.sink16_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.sink16_endofpacket   (rsp_xbar_demux_016_src0_endofpacket),   //          .endofpacket
		.sink17_ready         (rsp_xbar_demux_017_src0_ready),         //    sink17.ready
		.sink17_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.sink17_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.sink17_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.sink17_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.sink17_endofpacket   (rsp_xbar_demux_017_src0_endofpacket),   //          .endofpacket
		.sink18_ready         (rsp_xbar_demux_018_src0_ready),         //    sink18.ready
		.sink18_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.sink18_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.sink18_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.sink18_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.sink18_endofpacket   (rsp_xbar_demux_018_src0_endofpacket),   //          .endofpacket
		.sink19_ready         (rsp_xbar_demux_019_src0_ready),         //    sink19.ready
		.sink19_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.sink19_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.sink19_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.sink19_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.sink19_endofpacket   (rsp_xbar_demux_019_src0_endofpacket),   //          .endofpacket
		.sink20_ready         (rsp_xbar_demux_020_src0_ready),         //    sink20.ready
		.sink20_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.sink20_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.sink20_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.sink20_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.sink20_endofpacket   (rsp_xbar_demux_020_src0_endofpacket),   //          .endofpacket
		.sink21_ready         (rsp_xbar_demux_021_src0_ready),         //    sink21.ready
		.sink21_valid         (rsp_xbar_demux_021_src0_valid),         //          .valid
		.sink21_channel       (rsp_xbar_demux_021_src0_channel),       //          .channel
		.sink21_data          (rsp_xbar_demux_021_src0_data),          //          .data
		.sink21_startofpacket (rsp_xbar_demux_021_src0_startofpacket), //          .startofpacket
		.sink21_endofpacket   (rsp_xbar_demux_021_src0_endofpacket),   //          .endofpacket
		.sink22_ready         (rsp_xbar_demux_022_src0_ready),         //    sink22.ready
		.sink22_valid         (rsp_xbar_demux_022_src0_valid),         //          .valid
		.sink22_channel       (rsp_xbar_demux_022_src0_channel),       //          .channel
		.sink22_data          (rsp_xbar_demux_022_src0_data),          //          .data
		.sink22_startofpacket (rsp_xbar_demux_022_src0_startofpacket), //          .startofpacket
		.sink22_endofpacket   (rsp_xbar_demux_022_src0_endofpacket),   //          .endofpacket
		.sink23_ready         (rsp_xbar_demux_023_src0_ready),         //    sink23.ready
		.sink23_valid         (rsp_xbar_demux_023_src0_valid),         //          .valid
		.sink23_channel       (rsp_xbar_demux_023_src0_channel),       //          .channel
		.sink23_data          (rsp_xbar_demux_023_src0_data),          //          .data
		.sink23_startofpacket (rsp_xbar_demux_023_src0_startofpacket), //          .startofpacket
		.sink23_endofpacket   (rsp_xbar_demux_023_src0_endofpacket),   //          .endofpacket
		.sink24_ready         (rsp_xbar_demux_024_src0_ready),         //    sink24.ready
		.sink24_valid         (rsp_xbar_demux_024_src0_valid),         //          .valid
		.sink24_channel       (rsp_xbar_demux_024_src0_channel),       //          .channel
		.sink24_data          (rsp_xbar_demux_024_src0_data),          //          .data
		.sink24_startofpacket (rsp_xbar_demux_024_src0_startofpacket), //          .startofpacket
		.sink24_endofpacket   (rsp_xbar_demux_024_src0_endofpacket),   //          .endofpacket
		.sink25_ready         (rsp_xbar_demux_025_src0_ready),         //    sink25.ready
		.sink25_valid         (rsp_xbar_demux_025_src0_valid),         //          .valid
		.sink25_channel       (rsp_xbar_demux_025_src0_channel),       //          .channel
		.sink25_data          (rsp_xbar_demux_025_src0_data),          //          .data
		.sink25_startofpacket (rsp_xbar_demux_025_src0_startofpacket), //          .startofpacket
		.sink25_endofpacket   (rsp_xbar_demux_025_src0_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (61),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (70),
		.IN_PKT_BYTE_CNT_L             (68),
		.IN_PKT_TRANS_COMPRESSED_READ  (62),
		.IN_PKT_BURSTWRAP_H            (73),
		.IN_PKT_BURSTWRAP_L            (71),
		.IN_PKT_BURST_SIZE_H           (76),
		.IN_PKT_BURST_SIZE_L           (74),
		.IN_PKT_RESPONSE_STATUS_H      (102),
		.IN_PKT_RESPONSE_STATUS_L      (101),
		.IN_PKT_TRANS_EXCLUSIVE        (67),
		.IN_PKT_BURST_TYPE_H           (78),
		.IN_PKT_BURST_TYPE_L           (77),
		.IN_ST_DATA_W                  (103),
		.OUT_PKT_ADDR_H                (43),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (52),
		.OUT_PKT_BYTE_CNT_L            (50),
		.OUT_PKT_TRANS_COMPRESSED_READ (44),
		.OUT_PKT_BURST_SIZE_H          (58),
		.OUT_PKT_BURST_SIZE_L          (56),
		.OUT_PKT_RESPONSE_STATUS_H     (84),
		.OUT_PKT_RESPONSE_STATUS_L     (83),
		.OUT_PKT_TRANS_EXCLUSIVE       (49),
		.OUT_PKT_BURST_TYPE_H          (60),
		.OUT_PKT_BURST_TYPE_L          (59),
		.OUT_ST_DATA_W                 (85),
		.ST_CHANNEL_W                  (26),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter (
		.clk                  (altpll_0_c0_clk),                    //       clk.clk
		.reset                (rst_controller_001_reset_out_reset), // clk_reset.reset
		.in_valid             (cmd_xbar_mux_001_src_valid),         //      sink.valid
		.in_channel           (cmd_xbar_mux_001_src_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_mux_001_src_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_mux_001_src_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_mux_001_src_ready),         //          .ready
		.in_data              (cmd_xbar_mux_001_src_data),          //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_src_data),             //          .data
		.out_channel          (width_adapter_src_channel),          //          .channel
		.out_valid            (width_adapter_src_valid),            //          .valid
		.out_ready            (width_adapter_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                              // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (43),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (52),
		.IN_PKT_BYTE_CNT_L             (50),
		.IN_PKT_TRANS_COMPRESSED_READ  (44),
		.IN_PKT_BURSTWRAP_H            (55),
		.IN_PKT_BURSTWRAP_L            (53),
		.IN_PKT_BURST_SIZE_H           (58),
		.IN_PKT_BURST_SIZE_L           (56),
		.IN_PKT_RESPONSE_STATUS_H      (84),
		.IN_PKT_RESPONSE_STATUS_L      (83),
		.IN_PKT_TRANS_EXCLUSIVE        (49),
		.IN_PKT_BURST_TYPE_H           (60),
		.IN_PKT_BURST_TYPE_L           (59),
		.IN_ST_DATA_W                  (85),
		.OUT_PKT_ADDR_H                (61),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (70),
		.OUT_PKT_BYTE_CNT_L            (68),
		.OUT_PKT_TRANS_COMPRESSED_READ (62),
		.OUT_PKT_BURST_SIZE_H          (76),
		.OUT_PKT_BURST_SIZE_L          (74),
		.OUT_PKT_RESPONSE_STATUS_H     (102),
		.OUT_PKT_RESPONSE_STATUS_L     (101),
		.OUT_PKT_TRANS_EXCLUSIVE       (67),
		.OUT_PKT_BURST_TYPE_H          (78),
		.OUT_PKT_BURST_TYPE_L          (77),
		.OUT_ST_DATA_W                 (103),
		.ST_CHANNEL_W                  (26),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_001 (
		.clk                  (altpll_0_c0_clk),                     //       clk.clk
		.reset                (rst_controller_001_reset_out_reset),  // clk_reset.reset
		.in_valid             (id_router_001_src_valid),             //      sink.valid
		.in_channel           (id_router_001_src_channel),           //          .channel
		.in_startofpacket     (id_router_001_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_001_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_001_src_ready),             //          .ready
		.in_data              (id_router_001_src_data),              //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_001_src_data),          //          .data
		.out_channel          (width_adapter_001_src_channel),       //          .channel
		.out_valid            (width_adapter_001_src_valid),         //          .valid
		.out_ready            (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (26),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser (
		.in_clk            (altpll_0_c0_clk),                        //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),         //  in_clk_reset.reset
		.out_clk           (altpll_0_c2_clk),                        //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset),     // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src11_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src11_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src11_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src11_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src11_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src11_data),          //              .data
		.out_ready         (crosser_out_ready),                      //           out.ready
		.out_valid         (crosser_out_valid),                      //              .valid
		.out_startofpacket (crosser_out_startofpacket),              //              .startofpacket
		.out_endofpacket   (crosser_out_endofpacket),                //              .endofpacket
		.out_channel       (crosser_out_channel),                    //              .channel
		.out_data          (crosser_out_data),                       //              .data
		.in_empty          (1'b0),                                   //   (terminated)
		.in_error          (1'b0),                                   //   (terminated)
		.out_empty         (),                                       //   (terminated)
		.out_error         ()                                        //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (26),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_001 (
		.in_clk            (altpll_0_c2_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_0_c0_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_011_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_011_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_011_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_011_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_011_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_011_src0_data),          //              .data
		.out_ready         (crosser_001_out_ready),                 //           out.ready
		.out_valid         (crosser_001_out_valid),                 //              .valid
		.out_startofpacket (crosser_001_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_001_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_001_out_channel),               //              .channel
		.out_data          (crosser_001_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	NIOS_Sys_irq_mapper irq_mapper (
		.clk           (altpll_0_c0_clk),                //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.sender_irq    (nios2_qsys_0_d_irq_irq)          //    sender.irq
	);

endmodule
